`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company:
// Engineer:
//
// Create Date: 03/04/2024 09:10:17 AM
// Design Name:
// Module Name: EchoStateNetwork
// Project Name:
// Target Devices:
// Tool Versions:
// Description:
//
// Dependencies:
//
// Revision:
// Revision 0.01 - File Created
// Additional Comments:
//
//////////////////////////////////////////////////////////////////////////////////

module ESN_Generator_V2(
    input clk,
    input signed [7:0] input_data,     // Q2.6 format
    output wire signed [31:0] output_data   // Q2.6 format
);
parameter num_reservoir_neurons = 200;

// Reservoir layer
reg signed [15:0] a_scaled = 16'd-16384;
reg signed [15:0] b_scaled = 16'd16384;
reg signed [15:0] c_scaled = 16'd-19248;
reg signed [15:0] d_scaled = 16'd19248;
reg signed [31:0] reservoir_state [0: num_reservoir_neurons-1]; // Q4.12 format
initial begin
reservoir_state[0] = -32'sd84;
reservoir_state[1] = -32'sd80;
reservoir_state[2] = -32'sd124;
reservoir_state[3] = -32'sd55;
reservoir_state[4] = 32'sd121;
reservoir_state[5] = 32'sd112;
reservoir_state[6] = 32'sd94;
reservoir_state[7] = 32'sd115;
reservoir_state[8] = 32'sd116;
reservoir_state[9] = -32'sd115;
reservoir_state[10] = 32'sd101;
reservoir_state[11] = -32'sd58;
reservoir_state[12] = -32'sd77;
reservoir_state[13] = -32'sd119;
reservoir_state[14] = -32'sd101;
reservoir_state[15] = 32'sd61;
reservoir_state[16] = 32'sd71;
reservoir_state[17] = 32'sd54;
reservoir_state[18] = 32'sd116;
reservoir_state[19] = -32'sd95;
reservoir_state[20] = -32'sd101;
reservoir_state[21] = -32'sd122;
reservoir_state[22] = -32'sd113;
reservoir_state[23] = -32'sd101;
reservoir_state[24] = -32'sd121;
reservoir_state[25] = 32'sd31;
reservoir_state[26] = 32'sd124;
reservoir_state[27] = -32'sd5;
reservoir_state[28] = -32'sd126;
reservoir_state[29] = 32'sd101;
reservoir_state[30] = 32'sd70;
reservoir_state[31] = -32'sd6;
reservoir_state[32] = -32'sd94;
reservoir_state[33] = 32'sd124;
reservoir_state[34] = 32'sd84;
reservoir_state[35] = -32'sd124;
reservoir_state[36] = 32'sd105;
reservoir_state[37] = -32'sd69;
reservoir_state[38] = 32'sd89;
reservoir_state[39] = -32'sd33;
reservoir_state[40] = -32'sd65;
reservoir_state[41] = 32'sd109;
reservoir_state[42] = -32'sd126;
reservoir_state[43] = 32'sd76;
reservoir_state[44] = 32'sd81;
reservoir_state[45] = 32'sd111;
reservoir_state[46] = -32'sd84;
reservoir_state[47] = 32'sd62;
reservoir_state[48] = 32'sd111;
reservoir_state[49] = -32'sd105;
reservoir_state[50] = 32'sd120;
reservoir_state[51] = 32'sd115;
reservoir_state[52] = 32'sd90;
reservoir_state[53] = 32'sd38;
reservoir_state[54] = 32'sd127;
reservoir_state[55] = -32'sd126;
reservoir_state[56] = -32'sd43;
reservoir_state[57] = -32'sd86;
reservoir_state[58] = 32'sd122;
reservoir_state[59] = -32'sd29;
reservoir_state[60] = -32'sd110;
reservoir_state[61] = 32'sd14;
reservoir_state[62] = -32'sd89;
reservoir_state[63] = -32'sd107;
reservoir_state[64] = 32'sd1;
reservoir_state[65] = 32'sd117;
reservoir_state[66] = 32'sd124;
reservoir_state[67] = 32'sd108;
reservoir_state[68] = 32'sd115;
reservoir_state[69] = 32'sd108;
reservoir_state[70] = -32'sd82;
reservoir_state[71] = 32'sd60;
reservoir_state[72] = -32'sd40;
reservoir_state[73] = -32'sd118;
reservoir_state[74] = 32'sd72;
reservoir_state[75] = -32'sd107;
reservoir_state[76] = 32'sd67;
reservoir_state[77] = 32'sd117;
reservoir_state[78] = -32'sd121;
reservoir_state[79] = 32'sd104;
reservoir_state[80] = 32'sd77;
reservoir_state[81] = 32'sd119;
reservoir_state[82] = 32'sd112;
reservoir_state[83] = 32'sd83;
reservoir_state[84] = -32'sd125;
reservoir_state[85] = 32'sd92;
reservoir_state[86] = 32'sd9;
reservoir_state[87] = 32'sd91;
reservoir_state[88] = 32'sd114;
reservoir_state[89] = -32'sd123;
reservoir_state[90] = -32'sd90;
reservoir_state[91] = -32'sd9;
reservoir_state[92] = 32'sd127;
reservoir_state[93] = -32'sd77;
reservoir_state[94] = 32'sd105;
reservoir_state[95] = 32'sd46;
reservoir_state[96] = -32'sd62;
reservoir_state[97] = -32'sd106;
reservoir_state[98] = 32'sd87;
reservoir_state[99] = -32'sd104;
reservoir_state[100] = -32'sd82;
reservoir_state[101] = -32'sd88;
reservoir_state[102] = 32'sd126;
reservoir_state[103] = -32'sd64;
reservoir_state[104] = 32'sd11;
reservoir_state[105] = 32'sd116;
reservoir_state[106] = -32'sd126;
reservoir_state[107] = 32'sd87;
reservoir_state[108] = 32'sd96;
reservoir_state[109] = 32'sd80;
reservoir_state[110] = -32'sd116;
reservoir_state[111] = -32'sd80;
reservoir_state[112] = 32'sd119;
reservoir_state[113] = 32'sd115;
reservoir_state[114] = -32'sd45;
reservoir_state[115] = 32'sd38;
reservoir_state[116] = -32'sd24;
reservoir_state[117] = -32'sd111;
reservoir_state[118] = 32'sd114;
reservoir_state[119] = -32'sd111;
reservoir_state[120] = 32'sd103;
reservoir_state[121] = 32'sd51;
reservoir_state[122] = -32'sd82;
reservoir_state[123] = 32'sd58;
reservoir_state[124] = 32'sd23;
reservoir_state[125] = -32'sd61;
reservoir_state[126] = -32'sd119;
reservoir_state[127] = 32'sd10;
reservoir_state[128] = -32'sd117;
reservoir_state[129] = 32'sd112;
reservoir_state[130] = -32'sd34;
reservoir_state[131] = -32'sd100;
reservoir_state[132] = 32'sd82;
reservoir_state[133] = 32'sd127;
reservoir_state[134] = 32'sd32;
reservoir_state[135] = 32'sd93;
reservoir_state[136] = -32'sd110;
reservoir_state[137] = 32'sd79;
reservoir_state[138] = -32'sd20;
reservoir_state[139] = 32'sd52;
reservoir_state[140] = -32'sd71;
reservoir_state[141] = -32'sd124;
reservoir_state[142] = -32'sd10;
reservoir_state[143] = 32'sd119;
reservoir_state[144] = -32'sd105;
reservoir_state[145] = 32'sd14;
reservoir_state[146] = 32'sd122;
reservoir_state[147] = -32'sd46;
reservoir_state[148] = -32'sd121;
reservoir_state[149] = 32'sd100;
reservoir_state[150] = 32'sd71;
reservoir_state[151] = -32'sd99;
reservoir_state[152] = 32'sd104;
reservoir_state[153] = 32'sd73;
reservoir_state[154] = -32'sd104;
reservoir_state[155] = -32'sd127;
reservoir_state[156] = -32'sd111;
reservoir_state[157] = -32'sd93;
reservoir_state[158] = 32'sd26;
reservoir_state[159] = -32'sd87;
reservoir_state[160] = -32'sd7;
reservoir_state[161] = -32'sd92;
reservoir_state[162] = 32'sd89;
reservoir_state[163] = -32'sd16;
reservoir_state[164] = -32'sd43;
reservoir_state[165] = -32'sd107;
reservoir_state[166] = -32'sd122;
reservoir_state[167] = 32'sd127;
reservoir_state[168] = 32'sd111;
reservoir_state[169] = -32'sd123;
reservoir_state[170] = 32'sd8;
reservoir_state[171] = 32'sd126;
reservoir_state[172] = -32'sd123;
reservoir_state[173] = 32'sd16;
reservoir_state[174] = -32'sd127;
reservoir_state[175] = -32'sd116;
reservoir_state[176] = 32'sd65;
reservoir_state[177] = 32'sd126;
reservoir_state[178] = 32'sd112;
reservoir_state[179] = 32'sd118;
reservoir_state[180] = 32'sd71;
reservoir_state[181] = -32'sd106;
reservoir_state[182] = 32'sd23;
reservoir_state[183] = 32'sd60;
reservoir_state[184] = 32'sd127;
reservoir_state[185] = 32'sd104;
reservoir_state[186] = 32'sd107;
reservoir_state[187] = -32'sd85;
reservoir_state[188] = -32'sd108;
reservoir_state[189] = -32'sd68;
reservoir_state[190] = -32'sd82;
reservoir_state[191] = 32'sd98;
reservoir_state[192] = 32'sd114;
reservoir_state[193] = 32'sd119;
reservoir_state[194] = 32'sd110;
reservoir_state[195] = 32'sd57;
reservoir_state[196] = -32'sd78;
reservoir_state[197] = 32'sd19;
reservoir_state[198] = -32'sd128;
reservoir_state[199] = -32'sd92;
end

  // Scaling factors and zero point
  reg signed [31:0] scale = 32'b00000000000001011001011001000000;         // Q2.14 format

  reg signed [31:0] input_sum_parallel [0: num_reservoir_neurons-1];
  reg signed [31:0] reservoir_sum_parallel [0: num_reservoir_neurons-1];
  reg signed [31:0] output_sum;
  integer i,j,k,l,m;

  reg signed [31:0] reg_input [0: num_reservoir_neurons-1];
  reg signed [31:0] reg_reservoir [0: num_reservoir_neurons-1];
wire signed [31:0] shifted_state0_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state0_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state0_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state0_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state0_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state0_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state0_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state0_40_2 = reservoir_state[40] <<< 2;
wire signed [31:0] shifted_state0_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state0_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state0_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state0_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state0_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state0_47_4 = reservoir_state[47] <<< 4;
wire signed [31:0] shifted_state0_47_5 = reservoir_state[47] <<< 5;
wire signed [31:0] shifted_state0_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state0_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state0_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state0_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state0_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state0_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state0_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state0_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state0_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state0_87_3 = reservoir_state[87] <<< 3;
wire signed [31:0] shifted_state0_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state0_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state0_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state0_115_4 = reservoir_state[115] <<< 4;
wire signed [31:0] shifted_state0_115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state0_115_6 = reservoir_state[115] <<< 6;
wire signed [31:0] shifted_state0_115_7 = reservoir_state[115] <<< 7;
wire signed [31:0] shifted_state0_117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state0_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state0_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state0_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state0_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state0_117_5 = reservoir_state[117] <<< 5;
wire signed [31:0] shifted_state0_117_6 = reservoir_state[117] <<< 6;
wire signed [31:0] shifted_state0_117_7 = reservoir_state[117] <<< 7;
wire signed [31:0] shifted_state0_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state0_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state0_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state0_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state0_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state0_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state0_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state0_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state0_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state0_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state0_171_0 = reservoir_state[171] <<< 0;
wire signed [31:0] shifted_state0_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state0_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state0_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state0_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state0_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state0_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state0_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state0_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state0_176_2 = reservoir_state[176] <<< 2;
wire signed [31:0] shifted_state0_176_5 = reservoir_state[176] <<< 5;
wire signed [31:0] shifted_state0_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state0_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state0_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state0_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state0_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state0_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state0_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state0_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state0_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state0_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state0_196_3 = reservoir_state[196] <<< 3;
wire signed [31:0] shifted_state0_196_6 = reservoir_state[196] <<< 6;
wire signed [31:0] shifted_state1_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state1_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state1_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state1_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state1_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state1_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state1_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state1_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state1_12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state1_12_4 = reservoir_state[12] <<< 4;
wire signed [31:0] shifted_state1_14_0 = reservoir_state[14] <<< 0;
wire signed [31:0] shifted_state1_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state1_14_3 = reservoir_state[14] <<< 3;
wire signed [31:0] shifted_state1_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state1_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state1_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state1_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state1_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state1_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state1_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state1_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state1_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state1_57_3 = reservoir_state[57] <<< 3;
wire signed [31:0] shifted_state1_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state1_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state1_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state1_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state1_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state1_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state1_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state1_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state1_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state1_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state1_91_1 = reservoir_state[91] <<< 1;
wire signed [31:0] shifted_state1_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state1_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state1_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state1_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state1_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state1_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state1_93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state1_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state1_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state1_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state1_114_1 = reservoir_state[114] <<< 1;
wire signed [31:0] shifted_state1_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state1_119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state1_119_2 = reservoir_state[119] <<< 2;
wire signed [31:0] shifted_state1_119_3 = reservoir_state[119] <<< 3;
wire signed [31:0] shifted_state1_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state1_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state1_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state1_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state1_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state1_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state1_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state1_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state1_131_2 = reservoir_state[131] <<< 2;
wire signed [31:0] shifted_state1_131_4 = reservoir_state[131] <<< 4;
wire signed [31:0] shifted_state1_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state1_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state1_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state1_154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state1_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state1_154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state1_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state1_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state1_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state1_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state1_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state1_156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state1_156_6 = reservoir_state[156] <<< 6;
wire signed [31:0] shifted_state1_156_7 = reservoir_state[156] <<< 7;
wire signed [31:0] shifted_state1_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state1_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state1_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state1_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state1_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state1_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state1_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state1_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state1_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state1_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state2_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state2_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state2_17_4 = reservoir_state[17] <<< 4;
wire signed [31:0] shifted_state2_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state2_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state2_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state2_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state2_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state2_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state2_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state2_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state2_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state2_73_1 = reservoir_state[73] <<< 1;
wire signed [31:0] shifted_state2_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state2_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state2_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state2_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state2_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state2_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state2_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state2_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state2_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state2_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state2_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state2_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state2_140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state2_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state2_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state2_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state2_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state2_151_4 = reservoir_state[151] <<< 4;
wire signed [31:0] shifted_state2_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state2_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state2_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state2_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state2_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state2_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state2_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state2_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state2_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state2_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state2_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state2_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state2_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state2_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state2_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state2_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state3_15_1 = reservoir_state[15] <<< 1;
wire signed [31:0] shifted_state3_15_6 = reservoir_state[15] <<< 6;
wire signed [31:0] shifted_state3_15_7 = reservoir_state[15] <<< 7;
wire signed [31:0] shifted_state3_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state3_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state3_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state3_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state3_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state3_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state3_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state3_36_4 = reservoir_state[36] <<< 4;
wire signed [31:0] shifted_state3_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state3_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state3_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state3_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state3_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state3_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state3_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state3_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state3_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state3_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state3_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state3_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state3_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state3_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state3_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state3_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state3_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state3_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state3_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state3_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state3_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state3_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state3_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state3_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state3_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state3_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state3_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state3_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state3_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state3_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state3_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state3_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state3_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state3_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state3_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state3_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state3_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state3_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state3_149_5 = reservoir_state[149] <<< 5;
wire signed [31:0] shifted_state3_149_6 = reservoir_state[149] <<< 6;
wire signed [31:0] shifted_state3_149_7 = reservoir_state[149] <<< 7;
wire signed [31:0] shifted_state3_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state3_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state3_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state3_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state3_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state3_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state3_186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state3_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state3_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state3_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state3_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state3_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state3_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state3_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state4_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state4_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state4_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state4_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state4_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state4_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state4_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state4_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state4_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state4_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state4_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state4_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state4_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state4_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state4_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state4_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state4_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state4_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state4_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state4_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state4_58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state4_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state4_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state4_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state4_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state4_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state4_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state4_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state4_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state4_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state4_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state4_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state4_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state4_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state4_85_3 = reservoir_state[85] <<< 3;
wire signed [31:0] shifted_state4_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state4_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state4_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state4_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state4_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state4_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state4_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state4_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state4_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state4_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state4_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state4_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state4_119_3 = reservoir_state[119] <<< 3;
wire signed [31:0] shifted_state4_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state4_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state4_119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state4_119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state4_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state4_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state4_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state4_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state4_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state4_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state4_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state4_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state4_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state4_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state4_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state4_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state4_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state4_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state4_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state4_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state4_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state4_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state4_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state4_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state4_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state4_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state4_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state4_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state4_197_0 = reservoir_state[197] <<< 0;
wire signed [31:0] shifted_state4_197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state4_197_4 = reservoir_state[197] <<< 4;
wire signed [31:0] shifted_state4_197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state4_199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state4_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state4_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state4_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state4_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state4_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state5_12_0 = reservoir_state[12] <<< 0;
wire signed [31:0] shifted_state5_12_2 = reservoir_state[12] <<< 2;
wire signed [31:0] shifted_state5_12_4 = reservoir_state[12] <<< 4;
wire signed [31:0] shifted_state5_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state5_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state5_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state5_128_6 = reservoir_state[128] <<< 6;
wire signed [31:0] shifted_state5_128_7 = reservoir_state[128] <<< 7;
wire signed [31:0] shifted_state5_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state5_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state5_135_3 = reservoir_state[135] <<< 3;
wire signed [31:0] shifted_state5_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state5_143_0 = reservoir_state[143] <<< 0;
wire signed [31:0] shifted_state5_143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state5_143_2 = reservoir_state[143] <<< 2;
wire signed [31:0] shifted_state5_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state5_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state5_145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state5_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state5_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state5_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state5_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state5_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state5_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state5_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state5_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state5_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state5_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state5_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state5_162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state5_162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state5_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state5_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state5_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state5_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state5_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state5_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state5_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state5_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state5_199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state5_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state5_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state5_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state5_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state6_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state6_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state6_12_0 = reservoir_state[12] <<< 0;
wire signed [31:0] shifted_state6_12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state6_12_2 = reservoir_state[12] <<< 2;
wire signed [31:0] shifted_state6_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state6_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state6_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state6_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state6_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state6_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state6_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state6_64_4 = reservoir_state[64] <<< 4;
wire signed [31:0] shifted_state6_69_1 = reservoir_state[69] <<< 1;
wire signed [31:0] shifted_state6_69_2 = reservoir_state[69] <<< 2;
wire signed [31:0] shifted_state6_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state6_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state6_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state6_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state6_88_5 = reservoir_state[88] <<< 5;
wire signed [31:0] shifted_state6_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state6_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state6_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state6_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state6_112_3 = reservoir_state[112] <<< 3;
wire signed [31:0] shifted_state6_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state6_112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state6_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state6_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state6_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state6_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state6_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state6_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state6_147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state6_147_3 = reservoir_state[147] <<< 3;
wire signed [31:0] shifted_state6_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state6_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state6_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state6_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state6_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state6_158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state6_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state6_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state6_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state6_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state6_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state6_181_1 = reservoir_state[181] <<< 1;
wire signed [31:0] shifted_state6_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state6_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state6_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state6_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state6_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state6_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state6_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state6_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state6_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state6_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state6_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state6_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state7_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state7_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state7_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state7_16_3 = reservoir_state[16] <<< 3;
wire signed [31:0] shifted_state7_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state7_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state7_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state7_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state7_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state7_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state7_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state7_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state7_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state7_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state7_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state7_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state7_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state7_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state7_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state7_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state7_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state7_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state7_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state7_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state7_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state7_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state7_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state7_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state7_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state7_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state7_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state7_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state7_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state7_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state7_94_2 = reservoir_state[94] <<< 2;
wire signed [31:0] shifted_state7_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state7_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state7_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state7_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state7_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state7_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state7_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state7_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state7_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state7_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state7_128_2 = reservoir_state[128] <<< 2;
wire signed [31:0] shifted_state7_128_3 = reservoir_state[128] <<< 3;
wire signed [31:0] shifted_state7_128_5 = reservoir_state[128] <<< 5;
wire signed [31:0] shifted_state7_128_6 = reservoir_state[128] <<< 6;
wire signed [31:0] shifted_state7_128_7 = reservoir_state[128] <<< 7;
wire signed [31:0] shifted_state7_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state7_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state7_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state7_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state7_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state7_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state7_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state7_171_5 = reservoir_state[171] <<< 5;
wire signed [31:0] shifted_state7_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state7_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state7_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state7_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state7_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state7_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state8_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state8_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state8_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state8_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state8_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state8_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state8_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state8_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state8_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state8_36_1 = reservoir_state[36] <<< 1;
wire signed [31:0] shifted_state8_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state8_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state8_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state8_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state8_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state8_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state8_53_3 = reservoir_state[53] <<< 3;
wire signed [31:0] shifted_state8_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state8_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state8_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state8_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state8_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state8_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state8_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state8_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state8_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state8_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state8_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state8_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state8_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state8_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state8_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state8_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state8_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state8_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state8_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state8_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state8_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state8_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state8_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state8_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state8_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state8_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state8_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state8_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state8_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state8_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state8_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state8_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state8_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state8_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state8_114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state8_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state8_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state8_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state8_125_2 = reservoir_state[125] <<< 2;
wire signed [31:0] shifted_state8_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state8_125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state8_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state8_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state8_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state8_131_2 = reservoir_state[131] <<< 2;
wire signed [31:0] shifted_state8_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state8_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state8_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state8_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state8_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state8_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state8_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state8_149_2 = reservoir_state[149] <<< 2;
wire signed [31:0] shifted_state8_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state8_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state8_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state8_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state8_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state8_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state8_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state8_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state8_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state8_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state8_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state8_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state8_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state8_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state8_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state9_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state9_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state9_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state9_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state9_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state9_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state9_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state9_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state9_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state9_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state9_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state9_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state9_52_0 = reservoir_state[52] <<< 0;
wire signed [31:0] shifted_state9_52_1 = reservoir_state[52] <<< 1;
wire signed [31:0] shifted_state9_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state9_52_4 = reservoir_state[52] <<< 4;
wire signed [31:0] shifted_state9_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state9_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state9_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state9_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state9_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state9_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state9_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state9_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state9_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state9_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state9_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state9_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state9_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state9_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state9_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state9_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state9_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state9_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state9_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state9_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state9_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state9_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state9_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state9_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state9_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state9_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state9_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state9_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state9_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state9_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state9_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state9_137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state9_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state9_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state9_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state9_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state9_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state9_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state9_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state9_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state9_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state9_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state9_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state9_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state9_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state9_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state9_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state9_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state9_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state9_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state9_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state9_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state9_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state9_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state9_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state9_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state9_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state9_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state9_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state9_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state9_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state9_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state9_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state9_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state10_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state10_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state10_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state10_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state10_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state10_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state10_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state10_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state10_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state10_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state10_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state10_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state10_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state10_56_0 = reservoir_state[56] <<< 0;
wire signed [31:0] shifted_state10_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state10_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state10_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state10_73_3 = reservoir_state[73] <<< 3;
wire signed [31:0] shifted_state10_73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state10_73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state10_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state10_74_3 = reservoir_state[74] <<< 3;
wire signed [31:0] shifted_state10_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state10_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state10_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state10_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state10_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state10_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state10_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state10_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state10_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state10_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state10_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state10_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state10_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state10_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state10_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state10_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state10_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state10_131_2 = reservoir_state[131] <<< 2;
wire signed [31:0] shifted_state10_131_4 = reservoir_state[131] <<< 4;
wire signed [31:0] shifted_state10_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state10_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state10_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state10_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state10_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state10_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state10_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state10_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state10_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state10_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state10_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state10_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state10_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state10_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state10_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state10_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state10_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state10_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state10_176_0 = reservoir_state[176] <<< 0;
wire signed [31:0] shifted_state10_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state10_176_4 = reservoir_state[176] <<< 4;
wire signed [31:0] shifted_state10_176_5 = reservoir_state[176] <<< 5;
wire signed [31:0] shifted_state10_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state10_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state10_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state10_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state10_179_2 = reservoir_state[179] <<< 2;
wire signed [31:0] shifted_state10_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state10_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state10_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state10_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state10_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state10_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state10_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state10_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state10_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state10_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state10_185_0 = reservoir_state[185] <<< 0;
wire signed [31:0] shifted_state10_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state10_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state10_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state10_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state10_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state10_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state10_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state10_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state11_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state11_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state11_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state11_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state11_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state11_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state11_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state11_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state11_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state11_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state11_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state11_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state11_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state11_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state11_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state11_33_4 = reservoir_state[33] <<< 4;
wire signed [31:0] shifted_state11_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state11_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state11_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state11_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state11_34_2 = reservoir_state[34] <<< 2;
wire signed [31:0] shifted_state11_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state11_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state11_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state11_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state11_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state11_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state11_58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state11_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state11_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state11_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state11_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state11_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state11_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state11_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state11_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state11_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state11_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state11_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state11_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state11_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state11_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state11_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state11_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state11_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state11_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state11_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state11_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state11_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state11_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state11_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state11_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state11_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state11_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state11_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state11_135_4 = reservoir_state[135] <<< 4;
wire signed [31:0] shifted_state11_135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state11_135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state11_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state11_143_3 = reservoir_state[143] <<< 3;
wire signed [31:0] shifted_state11_143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state11_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state11_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state11_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state11_147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state11_147_5 = reservoir_state[147] <<< 5;
wire signed [31:0] shifted_state11_147_6 = reservoir_state[147] <<< 6;
wire signed [31:0] shifted_state11_147_7 = reservoir_state[147] <<< 7;
wire signed [31:0] shifted_state11_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state11_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state11_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state11_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state11_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state11_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state11_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state11_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state11_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state11_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state11_158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state11_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state12_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state12_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state12_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state12_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state12_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state12_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state12_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state12_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state12_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state12_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state12_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state12_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state12_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state12_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state12_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state12_54_4 = reservoir_state[54] <<< 4;
wire signed [31:0] shifted_state12_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state12_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state12_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state12_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state12_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state12_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state12_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state12_75_1 = reservoir_state[75] <<< 1;
wire signed [31:0] shifted_state12_75_2 = reservoir_state[75] <<< 2;
wire signed [31:0] shifted_state12_75_3 = reservoir_state[75] <<< 3;
wire signed [31:0] shifted_state12_75_5 = reservoir_state[75] <<< 5;
wire signed [31:0] shifted_state12_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state12_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state12_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state12_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state12_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state12_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state12_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state12_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state12_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state12_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state12_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state12_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state12_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state12_125_4 = reservoir_state[125] <<< 4;
wire signed [31:0] shifted_state12_125_5 = reservoir_state[125] <<< 5;
wire signed [31:0] shifted_state12_125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state12_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state12_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state12_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state12_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state12_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state12_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state12_144_0 = reservoir_state[144] <<< 0;
wire signed [31:0] shifted_state12_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state12_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state12_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state12_144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state12_144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state12_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state12_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state12_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state12_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state12_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state12_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state12_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state12_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state12_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state12_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state12_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state12_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state12_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state12_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state12_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state12_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state12_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state12_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state12_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state12_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state12_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state12_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state12_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state12_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state12_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state12_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state12_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state12_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state12_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state12_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state12_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state12_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state12_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state12_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state12_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state12_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state12_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state12_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state12_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state12_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state12_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state12_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state12_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state12_197_0 = reservoir_state[197] <<< 0;
wire signed [31:0] shifted_state12_197_2 = reservoir_state[197] <<< 2;
wire signed [31:0] shifted_state12_197_5 = reservoir_state[197] <<< 5;
wire signed [31:0] shifted_state12_199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state12_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state12_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state12_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state12_199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state12_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state12_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state12_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state13_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state13_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state13_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state13_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state13_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state13_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state13_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state13_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state13_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state13_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state13_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state13_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state13_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state13_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state13_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state13_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state13_27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state13_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state13_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state13_27_4 = reservoir_state[27] <<< 4;
wire signed [31:0] shifted_state13_27_5 = reservoir_state[27] <<< 5;
wire signed [31:0] shifted_state13_27_6 = reservoir_state[27] <<< 6;
wire signed [31:0] shifted_state13_27_7 = reservoir_state[27] <<< 7;
wire signed [31:0] shifted_state13_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state13_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state13_30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state13_30_4 = reservoir_state[30] <<< 4;
wire signed [31:0] shifted_state13_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state13_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state13_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state13_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state13_57_3 = reservoir_state[57] <<< 3;
wire signed [31:0] shifted_state13_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state13_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state13_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state13_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state13_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state13_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state13_79_5 = reservoir_state[79] <<< 5;
wire signed [31:0] shifted_state13_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state13_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state13_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state13_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state13_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state13_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state13_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state13_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state13_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state13_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state13_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state13_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state13_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state13_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state13_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state13_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state13_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state13_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state13_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state13_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state13_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state13_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state13_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state13_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state13_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state13_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state13_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state13_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state13_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state13_145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state13_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state13_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state13_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state13_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state13_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state13_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state13_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state13_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state14_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state14_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state14_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state14_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state14_30_5 = reservoir_state[30] <<< 5;
wire signed [31:0] shifted_state14_30_6 = reservoir_state[30] <<< 6;
wire signed [31:0] shifted_state14_30_7 = reservoir_state[30] <<< 7;
wire signed [31:0] shifted_state14_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state14_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state14_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state14_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state14_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state14_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state14_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state14_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state14_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state14_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state14_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state14_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state14_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state14_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state14_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state14_68_1 = reservoir_state[68] <<< 1;
wire signed [31:0] shifted_state14_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state14_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state14_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state14_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state14_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state14_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state14_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state14_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state14_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state14_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state14_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state14_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state14_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state14_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state14_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state14_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state14_120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state14_120_5 = reservoir_state[120] <<< 5;
wire signed [31:0] shifted_state14_120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state14_120_7 = reservoir_state[120] <<< 7;
wire signed [31:0] shifted_state14_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state14_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state14_183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state14_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state14_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state14_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state15_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state15_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state15_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state15_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state15_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state15_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state15_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state15_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state15_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state15_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state15_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state15_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state15_5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state15_5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state15_5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state15_5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state15_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state15_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state15_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state15_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state15_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state15_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state15_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state15_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state15_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state15_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state15_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state15_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state15_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state15_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state15_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state15_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state15_111_4 = reservoir_state[111] <<< 4;
wire signed [31:0] shifted_state15_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state15_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state15_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state15_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state15_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state15_114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state15_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state15_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state15_119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state15_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state15_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state15_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state15_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state15_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state15_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state15_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state15_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state15_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state15_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state15_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state15_154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state15_157_0 = reservoir_state[157] <<< 0;
wire signed [31:0] shifted_state15_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state15_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state15_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state15_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state15_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state15_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state15_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state15_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state15_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state15_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state15_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state15_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state15_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state15_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state15_197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state15_197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state15_197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state15_197_7 = reservoir_state[197] <<< 7;
wire signed [31:0] shifted_state15_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state16_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state16_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state16_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state16_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state16_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state16_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state16_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state16_36_1 = reservoir_state[36] <<< 1;
wire signed [31:0] shifted_state16_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state16_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state16_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state16_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state16_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state16_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state16_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state16_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state16_72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state16_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state16_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state16_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state16_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state16_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state16_79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state16_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state16_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state16_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state16_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state16_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state16_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state16_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state16_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state16_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state16_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state16_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state16_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state16_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state16_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state16_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state16_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state16_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state16_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state16_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state16_134_0 = reservoir_state[134] <<< 0;
wire signed [31:0] shifted_state16_134_4 = reservoir_state[134] <<< 4;
wire signed [31:0] shifted_state16_134_5 = reservoir_state[134] <<< 5;
wire signed [31:0] shifted_state16_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state16_134_7 = reservoir_state[134] <<< 7;
wire signed [31:0] shifted_state16_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state16_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state16_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state16_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state16_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state16_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state16_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state16_157_0 = reservoir_state[157] <<< 0;
wire signed [31:0] shifted_state16_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state16_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state16_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state16_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state16_159_1 = reservoir_state[159] <<< 1;
wire signed [31:0] shifted_state16_159_4 = reservoir_state[159] <<< 4;
wire signed [31:0] shifted_state16_159_5 = reservoir_state[159] <<< 5;
wire signed [31:0] shifted_state16_159_6 = reservoir_state[159] <<< 6;
wire signed [31:0] shifted_state16_159_7 = reservoir_state[159] <<< 7;
wire signed [31:0] shifted_state16_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state16_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state16_185_0 = reservoir_state[185] <<< 0;
wire signed [31:0] shifted_state16_185_2 = reservoir_state[185] <<< 2;
wire signed [31:0] shifted_state16_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state16_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state16_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state16_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state16_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state17_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state17_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state17_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state17_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state17_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state17_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state17_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state17_17_4 = reservoir_state[17] <<< 4;
wire signed [31:0] shifted_state17_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state17_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state17_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state17_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state17_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state17_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state17_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state17_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state17_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state17_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state17_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state17_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state17_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state17_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state17_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state17_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state17_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state17_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state17_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state17_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state17_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state17_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state17_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state17_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state17_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state17_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state17_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state17_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state17_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state17_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state17_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state17_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state17_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state17_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state17_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state17_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state17_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state17_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state17_93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state17_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state17_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state17_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state17_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state17_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state17_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state17_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state17_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state17_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state17_128_3 = reservoir_state[128] <<< 3;
wire signed [31:0] shifted_state17_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state17_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state17_140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state17_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state17_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state17_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state17_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state17_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state17_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state17_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state17_143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state17_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state17_160_1 = reservoir_state[160] <<< 1;
wire signed [31:0] shifted_state17_160_2 = reservoir_state[160] <<< 2;
wire signed [31:0] shifted_state17_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state17_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state17_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state17_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state17_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state17_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state17_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state17_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state17_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state17_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state17_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state17_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state17_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state17_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state17_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state17_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state17_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state17_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state17_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state17_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state17_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state17_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state17_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state17_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state17_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state17_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state18_3_1 = reservoir_state[3] <<< 1;
wire signed [31:0] shifted_state18_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state18_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state18_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state18_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state18_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state18_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state18_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state18_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state18_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state18_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state18_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state18_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state18_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state18_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state18_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state18_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state18_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state18_27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state18_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state18_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state18_27_5 = reservoir_state[27] <<< 5;
wire signed [31:0] shifted_state18_27_6 = reservoir_state[27] <<< 6;
wire signed [31:0] shifted_state18_27_7 = reservoir_state[27] <<< 7;
wire signed [31:0] shifted_state18_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state18_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state18_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state18_67_3 = reservoir_state[67] <<< 3;
wire signed [31:0] shifted_state18_67_4 = reservoir_state[67] <<< 4;
wire signed [31:0] shifted_state18_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state18_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state18_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state18_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state18_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state18_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state18_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state18_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state18_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state18_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state18_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state18_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state18_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state18_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state18_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state18_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state18_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state18_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state18_113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state18_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state18_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state18_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state18_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state18_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state18_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state18_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state18_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state18_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state18_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state18_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state18_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state18_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state18_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state18_135_3 = reservoir_state[135] <<< 3;
wire signed [31:0] shifted_state18_135_4 = reservoir_state[135] <<< 4;
wire signed [31:0] shifted_state18_135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state18_135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state18_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state18_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state18_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state18_143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state18_143_2 = reservoir_state[143] <<< 2;
wire signed [31:0] shifted_state18_143_3 = reservoir_state[143] <<< 3;
wire signed [31:0] shifted_state18_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state18_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state18_151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state18_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state18_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state18_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state18_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state18_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state18_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state18_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state18_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state18_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state18_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state18_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state18_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state18_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state18_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state18_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state18_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state18_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state18_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state18_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state18_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state18_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state18_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state18_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state18_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state18_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state18_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state18_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state18_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state18_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state18_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state18_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state18_196_0 = reservoir_state[196] <<< 0;
wire signed [31:0] shifted_state18_196_1 = reservoir_state[196] <<< 1;
wire signed [31:0] shifted_state18_196_2 = reservoir_state[196] <<< 2;
wire signed [31:0] shifted_state18_196_4 = reservoir_state[196] <<< 4;
wire signed [31:0] shifted_state18_196_5 = reservoir_state[196] <<< 5;
wire signed [31:0] shifted_state18_196_6 = reservoir_state[196] <<< 6;
wire signed [31:0] shifted_state18_196_7 = reservoir_state[196] <<< 7;
wire signed [31:0] shifted_state19_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state19_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state19_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state19_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state19_27_5 = reservoir_state[27] <<< 5;
wire signed [31:0] shifted_state19_27_6 = reservoir_state[27] <<< 6;
wire signed [31:0] shifted_state19_27_7 = reservoir_state[27] <<< 7;
wire signed [31:0] shifted_state19_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state19_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state19_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state19_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state19_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state19_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state19_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state19_67_1 = reservoir_state[67] <<< 1;
wire signed [31:0] shifted_state19_67_4 = reservoir_state[67] <<< 4;
wire signed [31:0] shifted_state19_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state19_67_6 = reservoir_state[67] <<< 6;
wire signed [31:0] shifted_state19_67_7 = reservoir_state[67] <<< 7;
wire signed [31:0] shifted_state19_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state19_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state19_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state19_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state19_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state19_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state19_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state19_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state19_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state19_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state19_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state19_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state19_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state19_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state19_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state19_84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state19_84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state19_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state19_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state19_101_2 = reservoir_state[101] <<< 2;
wire signed [31:0] shifted_state19_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state19_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state19_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state19_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state19_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state19_110_0 = reservoir_state[110] <<< 0;
wire signed [31:0] shifted_state19_110_1 = reservoir_state[110] <<< 1;
wire signed [31:0] shifted_state19_110_2 = reservoir_state[110] <<< 2;
wire signed [31:0] shifted_state19_110_4 = reservoir_state[110] <<< 4;
wire signed [31:0] shifted_state19_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state19_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state19_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state19_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state19_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state19_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state19_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state19_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state19_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state19_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state19_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state19_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state19_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state19_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state19_140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state19_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state19_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state19_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state19_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state19_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state19_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state19_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state19_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state19_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state19_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state19_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state19_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state19_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state19_176_2 = reservoir_state[176] <<< 2;
wire signed [31:0] shifted_state19_176_4 = reservoir_state[176] <<< 4;
wire signed [31:0] shifted_state19_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state19_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state19_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state19_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state19_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state19_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state19_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state19_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state19_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state20_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state20_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state20_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state20_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state20_8_1 = reservoir_state[8] <<< 1;
wire signed [31:0] shifted_state20_8_3 = reservoir_state[8] <<< 3;
wire signed [31:0] shifted_state20_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state20_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state20_16_3 = reservoir_state[16] <<< 3;
wire signed [31:0] shifted_state20_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state20_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state20_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state20_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state20_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state20_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state20_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state20_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state20_27_0 = reservoir_state[27] <<< 0;
wire signed [31:0] shifted_state20_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state20_27_4 = reservoir_state[27] <<< 4;
wire signed [31:0] shifted_state20_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state20_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state20_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state20_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state20_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state20_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state20_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state20_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state20_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state20_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state20_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state20_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state20_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state20_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state20_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state20_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state20_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state20_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state20_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state20_158_0 = reservoir_state[158] <<< 0;
wire signed [31:0] shifted_state20_158_3 = reservoir_state[158] <<< 3;
wire signed [31:0] shifted_state20_160_1 = reservoir_state[160] <<< 1;
wire signed [31:0] shifted_state20_160_2 = reservoir_state[160] <<< 2;
wire signed [31:0] shifted_state20_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state20_169_2 = reservoir_state[169] <<< 2;
wire signed [31:0] shifted_state20_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state20_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state20_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state20_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state20_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state20_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state20_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state20_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state21_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state21_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state21_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state21_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state21_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state21_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state21_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state21_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state21_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state21_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state21_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state21_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state21_27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state21_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state21_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state21_27_4 = reservoir_state[27] <<< 4;
wire signed [31:0] shifted_state21_27_5 = reservoir_state[27] <<< 5;
wire signed [31:0] shifted_state21_27_6 = reservoir_state[27] <<< 6;
wire signed [31:0] shifted_state21_27_7 = reservoir_state[27] <<< 7;
wire signed [31:0] shifted_state21_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state21_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state21_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state21_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state21_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state21_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state21_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state21_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state21_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state21_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state21_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state21_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state21_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state21_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state21_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state21_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state21_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state21_75_1 = reservoir_state[75] <<< 1;
wire signed [31:0] shifted_state21_75_3 = reservoir_state[75] <<< 3;
wire signed [31:0] shifted_state21_75_4 = reservoir_state[75] <<< 4;
wire signed [31:0] shifted_state21_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state21_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state21_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state21_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state21_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state21_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state21_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state21_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state21_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state21_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state21_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state21_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state21_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state21_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state21_113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state21_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state21_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state21_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state21_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state21_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state21_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state21_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state21_124_2 = reservoir_state[124] <<< 2;
wire signed [31:0] shifted_state21_124_3 = reservoir_state[124] <<< 3;
wire signed [31:0] shifted_state21_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state21_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state21_124_6 = reservoir_state[124] <<< 6;
wire signed [31:0] shifted_state21_124_7 = reservoir_state[124] <<< 7;
wire signed [31:0] shifted_state21_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state21_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state21_134_5 = reservoir_state[134] <<< 5;
wire signed [31:0] shifted_state21_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state21_134_7 = reservoir_state[134] <<< 7;
wire signed [31:0] shifted_state21_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state21_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state21_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state21_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state21_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state21_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state21_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state21_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state21_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state21_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state21_158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state21_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state21_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state21_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state21_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state21_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state21_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state21_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state21_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state21_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state21_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state21_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state21_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state21_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state21_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state21_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state22_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state22_16_3 = reservoir_state[16] <<< 3;
wire signed [31:0] shifted_state22_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state22_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state22_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state22_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state22_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state22_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state22_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state22_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state22_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state22_30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state22_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state22_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state22_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state22_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state22_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state22_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state22_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state22_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state22_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state22_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state22_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state22_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state22_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state22_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state22_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state22_75_1 = reservoir_state[75] <<< 1;
wire signed [31:0] shifted_state22_75_2 = reservoir_state[75] <<< 2;
wire signed [31:0] shifted_state22_75_5 = reservoir_state[75] <<< 5;
wire signed [31:0] shifted_state22_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state22_92_1 = reservoir_state[92] <<< 1;
wire signed [31:0] shifted_state22_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state22_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state22_92_6 = reservoir_state[92] <<< 6;
wire signed [31:0] shifted_state22_92_7 = reservoir_state[92] <<< 7;
wire signed [31:0] shifted_state22_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state22_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state22_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state22_93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state22_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state22_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state22_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state22_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state22_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state22_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state22_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state22_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state22_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state22_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state22_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state22_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state22_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state22_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state22_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state22_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state22_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state22_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state22_167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state22_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state22_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state22_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state22_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state22_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state22_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state22_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state22_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state22_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state22_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state22_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state22_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state22_197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state22_199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state22_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state22_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state22_199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state22_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state22_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state22_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state23_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state23_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state23_9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state23_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state23_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state23_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state23_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state23_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state23_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state23_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state23_47_5 = reservoir_state[47] <<< 5;
wire signed [31:0] shifted_state23_56_0 = reservoir_state[56] <<< 0;
wire signed [31:0] shifted_state23_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state23_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state23_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state23_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state23_67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state23_67_1 = reservoir_state[67] <<< 1;
wire signed [31:0] shifted_state23_67_4 = reservoir_state[67] <<< 4;
wire signed [31:0] shifted_state23_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state23_67_6 = reservoir_state[67] <<< 6;
wire signed [31:0] shifted_state23_67_7 = reservoir_state[67] <<< 7;
wire signed [31:0] shifted_state23_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state23_88_5 = reservoir_state[88] <<< 5;
wire signed [31:0] shifted_state23_88_6 = reservoir_state[88] <<< 6;
wire signed [31:0] shifted_state23_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state23_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state23_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state23_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state23_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state23_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state23_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state23_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state23_101_2 = reservoir_state[101] <<< 2;
wire signed [31:0] shifted_state23_101_3 = reservoir_state[101] <<< 3;
wire signed [31:0] shifted_state23_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state23_102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state23_102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state23_102_7 = reservoir_state[102] <<< 7;
wire signed [31:0] shifted_state23_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state23_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state23_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state23_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state23_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state23_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state23_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state23_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state23_119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state23_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state23_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state23_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state23_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state23_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state23_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state23_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state23_140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state23_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state23_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state23_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state23_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state23_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state23_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state23_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state23_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state23_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state23_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state23_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state23_167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state23_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state23_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state23_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state23_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state23_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state23_181_3 = reservoir_state[181] <<< 3;
wire signed [31:0] shifted_state23_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state23_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state23_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state23_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state23_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state23_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state23_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state23_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state23_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state23_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state23_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state23_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state24_1_1 = reservoir_state[1] <<< 1;
wire signed [31:0] shifted_state24_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state24_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state24_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state24_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state24_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state24_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state24_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state24_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state24_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state24_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state24_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state24_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state24_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state24_9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state24_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state24_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state24_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state24_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state24_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state24_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state24_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state24_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state24_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state24_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state24_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state24_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state24_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state24_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state24_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state24_29_2 = reservoir_state[29] <<< 2;
wire signed [31:0] shifted_state24_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state24_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state24_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state24_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state24_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state24_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state24_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state24_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state24_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state24_49_1 = reservoir_state[49] <<< 1;
wire signed [31:0] shifted_state24_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state24_49_3 = reservoir_state[49] <<< 3;
wire signed [31:0] shifted_state24_49_4 = reservoir_state[49] <<< 4;
wire signed [31:0] shifted_state24_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state24_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state24_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state24_69_1 = reservoir_state[69] <<< 1;
wire signed [31:0] shifted_state24_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state24_69_5 = reservoir_state[69] <<< 5;
wire signed [31:0] shifted_state24_69_6 = reservoir_state[69] <<< 6;
wire signed [31:0] shifted_state24_69_7 = reservoir_state[69] <<< 7;
wire signed [31:0] shifted_state24_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state24_87_2 = reservoir_state[87] <<< 2;
wire signed [31:0] shifted_state24_87_3 = reservoir_state[87] <<< 3;
wire signed [31:0] shifted_state24_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state24_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state24_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state24_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state24_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state24_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state24_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state24_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state24_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state24_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state24_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state24_102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state24_102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state24_102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state24_102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state24_102_7 = reservoir_state[102] <<< 7;
wire signed [31:0] shifted_state24_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state24_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state24_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state24_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state24_131_2 = reservoir_state[131] <<< 2;
wire signed [31:0] shifted_state24_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state24_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state24_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state24_154_0 = reservoir_state[154] <<< 0;
wire signed [31:0] shifted_state24_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state24_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state24_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state24_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state24_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state24_169_2 = reservoir_state[169] <<< 2;
wire signed [31:0] shifted_state24_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state24_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state24_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state24_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state24_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state24_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state24_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state24_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state24_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state24_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state24_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state25_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state25_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state25_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state25_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state25_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state25_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state25_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state25_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state25_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state25_19_1 = reservoir_state[19] <<< 1;
wire signed [31:0] shifted_state25_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state25_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state25_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state25_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state25_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state25_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state25_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state25_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state25_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state25_50_4 = reservoir_state[50] <<< 4;
wire signed [31:0] shifted_state25_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state25_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state25_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state25_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state25_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state25_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state25_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state25_53_1 = reservoir_state[53] <<< 1;
wire signed [31:0] shifted_state25_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state25_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state25_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state25_75_1 = reservoir_state[75] <<< 1;
wire signed [31:0] shifted_state25_75_2 = reservoir_state[75] <<< 2;
wire signed [31:0] shifted_state25_75_4 = reservoir_state[75] <<< 4;
wire signed [31:0] shifted_state25_75_5 = reservoir_state[75] <<< 5;
wire signed [31:0] shifted_state25_75_6 = reservoir_state[75] <<< 6;
wire signed [31:0] shifted_state25_75_7 = reservoir_state[75] <<< 7;
wire signed [31:0] shifted_state25_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state25_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state25_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state25_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state25_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state25_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state25_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state25_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state25_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state25_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state25_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state25_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state25_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state25_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state25_122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state25_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state25_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state25_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state25_153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state25_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state25_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state25_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state25_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state25_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state25_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state25_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state25_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state25_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state25_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state25_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state25_185_0 = reservoir_state[185] <<< 0;
wire signed [31:0] shifted_state25_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state25_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state25_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state25_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state25_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state25_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state25_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state25_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state25_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state25_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state25_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state25_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state25_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state26_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state26_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state26_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state26_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state26_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state26_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state26_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state26_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state26_18_3 = reservoir_state[18] <<< 3;
wire signed [31:0] shifted_state26_27_0 = reservoir_state[27] <<< 0;
wire signed [31:0] shifted_state26_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state26_27_4 = reservoir_state[27] <<< 4;
wire signed [31:0] shifted_state26_27_5 = reservoir_state[27] <<< 5;
wire signed [31:0] shifted_state26_27_6 = reservoir_state[27] <<< 6;
wire signed [31:0] shifted_state26_27_7 = reservoir_state[27] <<< 7;
wire signed [31:0] shifted_state26_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state26_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state26_30_4 = reservoir_state[30] <<< 4;
wire signed [31:0] shifted_state26_30_6 = reservoir_state[30] <<< 6;
wire signed [31:0] shifted_state26_30_7 = reservoir_state[30] <<< 7;
wire signed [31:0] shifted_state26_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state26_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state26_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state26_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state26_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state26_54_4 = reservoir_state[54] <<< 4;
wire signed [31:0] shifted_state26_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state26_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state26_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state26_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state26_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state26_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state26_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state26_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state26_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state26_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state26_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state26_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state26_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state26_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state26_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state26_117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state26_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state26_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state26_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state26_117_6 = reservoir_state[117] <<< 6;
wire signed [31:0] shifted_state26_117_7 = reservoir_state[117] <<< 7;
wire signed [31:0] shifted_state26_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state26_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state26_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state26_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state26_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state26_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state26_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state26_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state26_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state26_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state26_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state27_2_0 = reservoir_state[2] <<< 0;
wire signed [31:0] shifted_state27_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state27_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state27_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state27_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state27_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state27_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state27_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state27_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state27_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state27_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state27_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state27_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state27_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state27_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state27_27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state27_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state27_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state27_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state27_65_2 = reservoir_state[65] <<< 2;
wire signed [31:0] shifted_state27_65_3 = reservoir_state[65] <<< 3;
wire signed [31:0] shifted_state27_65_5 = reservoir_state[65] <<< 5;
wire signed [31:0] shifted_state27_65_6 = reservoir_state[65] <<< 6;
wire signed [31:0] shifted_state27_65_7 = reservoir_state[65] <<< 7;
wire signed [31:0] shifted_state27_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state27_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state27_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state27_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state27_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state27_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state27_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state27_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state27_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state27_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state27_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state27_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state27_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state27_114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state27_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state27_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state27_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state27_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state27_117_5 = reservoir_state[117] <<< 5;
wire signed [31:0] shifted_state27_117_6 = reservoir_state[117] <<< 6;
wire signed [31:0] shifted_state27_117_7 = reservoir_state[117] <<< 7;
wire signed [31:0] shifted_state27_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state27_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state27_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state27_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state27_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state27_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state27_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state27_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state27_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state27_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state27_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state27_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state27_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state27_148_4 = reservoir_state[148] <<< 4;
wire signed [31:0] shifted_state27_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state27_148_6 = reservoir_state[148] <<< 6;
wire signed [31:0] shifted_state27_148_7 = reservoir_state[148] <<< 7;
wire signed [31:0] shifted_state27_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state27_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state27_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state27_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state27_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state27_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state27_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state27_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state27_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state27_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state27_176_3 = reservoir_state[176] <<< 3;
wire signed [31:0] shifted_state27_176_4 = reservoir_state[176] <<< 4;
wire signed [31:0] shifted_state27_176_5 = reservoir_state[176] <<< 5;
wire signed [31:0] shifted_state27_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state27_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state27_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state27_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state27_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state27_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state27_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state27_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state27_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state27_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state27_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state27_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state28_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state28_1_1 = reservoir_state[1] <<< 1;
wire signed [31:0] shifted_state28_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state28_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state28_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state28_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state28_2_0 = reservoir_state[2] <<< 0;
wire signed [31:0] shifted_state28_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state28_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state28_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state28_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state28_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state28_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state28_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state28_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state28_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state28_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state28_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state28_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state28_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state28_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state28_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state28_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state28_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state28_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state28_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state28_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state28_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state28_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state28_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state28_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state28_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state28_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state28_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state28_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state28_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state28_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state28_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state28_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state28_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state28_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state28_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state28_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state28_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state28_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state28_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state28_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state28_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state28_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state28_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state28_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state28_79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state28_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state28_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state28_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state28_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state28_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state28_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state28_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state28_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state28_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state28_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state28_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state28_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state28_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state28_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state28_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state28_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state28_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state28_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state28_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state28_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state28_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state28_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state28_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state28_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state28_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state28_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state28_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state28_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state28_140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state28_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state28_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state28_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state28_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state28_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state28_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state28_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state28_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state28_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state28_144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state28_144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state28_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state28_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state28_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state28_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state28_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state28_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state28_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state28_186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state28_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state28_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state28_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state28_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state28_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state28_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state28_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state28_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state28_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state28_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state28_189_6 = reservoir_state[189] <<< 6;
wire signed [31:0] shifted_state28_189_7 = reservoir_state[189] <<< 7;
wire signed [31:0] shifted_state28_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state28_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state28_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state28_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state28_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state28_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state28_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state29_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state29_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state29_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state29_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state29_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state29_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state29_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state29_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state29_14_3 = reservoir_state[14] <<< 3;
wire signed [31:0] shifted_state29_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state29_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state29_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state29_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state29_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state29_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state29_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state29_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state29_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state29_18_3 = reservoir_state[18] <<< 3;
wire signed [31:0] shifted_state29_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state29_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state29_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state29_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state29_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state29_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state29_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state29_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state29_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state29_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state29_49_1 = reservoir_state[49] <<< 1;
wire signed [31:0] shifted_state29_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state29_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state29_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state29_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state29_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state29_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state29_60_4 = reservoir_state[60] <<< 4;
wire signed [31:0] shifted_state29_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state29_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state29_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state29_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state29_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state29_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state29_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state29_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state29_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state29_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state29_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state29_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state29_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state29_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state29_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state29_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state29_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state29_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state29_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state29_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state29_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state29_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state29_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state29_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state29_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state29_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state29_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state29_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state29_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state29_171_0 = reservoir_state[171] <<< 0;
wire signed [31:0] shifted_state29_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state29_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state29_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state29_171_5 = reservoir_state[171] <<< 5;
wire signed [31:0] shifted_state29_171_6 = reservoir_state[171] <<< 6;
wire signed [31:0] shifted_state29_171_7 = reservoir_state[171] <<< 7;
wire signed [31:0] shifted_state29_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state29_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state29_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state29_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state29_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state29_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state29_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state29_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state29_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state29_183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state29_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state29_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state29_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state29_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state29_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state29_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state29_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state29_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state29_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state29_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state29_196_1 = reservoir_state[196] <<< 1;
wire signed [31:0] shifted_state29_196_4 = reservoir_state[196] <<< 4;
wire signed [31:0] shifted_state29_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state29_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state29_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state29_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state30_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state30_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state30_8_3 = reservoir_state[8] <<< 3;
wire signed [31:0] shifted_state30_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state30_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state30_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state30_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state30_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state30_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state30_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state30_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state30_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state30_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state30_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state30_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state30_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state30_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state30_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state30_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state30_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state30_64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state30_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state30_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state30_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state30_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state30_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state30_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state30_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state30_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state30_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state30_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state30_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state30_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state30_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state30_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state30_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state30_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state30_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state30_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state30_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state30_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state30_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state30_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state30_117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state30_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state30_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state30_117_5 = reservoir_state[117] <<< 5;
wire signed [31:0] shifted_state30_117_6 = reservoir_state[117] <<< 6;
wire signed [31:0] shifted_state30_117_7 = reservoir_state[117] <<< 7;
wire signed [31:0] shifted_state30_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state30_120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state30_120_5 = reservoir_state[120] <<< 5;
wire signed [31:0] shifted_state30_120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state30_120_7 = reservoir_state[120] <<< 7;
wire signed [31:0] shifted_state30_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state30_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state30_142_0 = reservoir_state[142] <<< 0;
wire signed [31:0] shifted_state30_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state30_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state30_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state30_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state30_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state30_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state30_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state30_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state30_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state30_151_4 = reservoir_state[151] <<< 4;
wire signed [31:0] shifted_state30_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state30_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state30_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state30_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state30_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state30_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state30_156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state30_156_6 = reservoir_state[156] <<< 6;
wire signed [31:0] shifted_state30_156_7 = reservoir_state[156] <<< 7;
wire signed [31:0] shifted_state30_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state30_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state30_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state30_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state30_169_2 = reservoir_state[169] <<< 2;
wire signed [31:0] shifted_state30_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state30_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state30_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state30_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state30_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state30_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state30_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state30_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state30_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state30_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state30_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state30_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state30_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state30_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state30_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state30_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state31_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state31_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state31_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state31_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state31_52_0 = reservoir_state[52] <<< 0;
wire signed [31:0] shifted_state31_52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state31_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state31_52_6 = reservoir_state[52] <<< 6;
wire signed [31:0] shifted_state31_56_0 = reservoir_state[56] <<< 0;
wire signed [31:0] shifted_state31_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state31_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state31_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state31_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state31_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state31_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state31_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state31_58_2 = reservoir_state[58] <<< 2;
wire signed [31:0] shifted_state31_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state31_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state31_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state31_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state31_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state31_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state31_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state31_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state31_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state31_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state31_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state31_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state31_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state31_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state31_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state31_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state31_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state31_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state31_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state31_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state31_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state31_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state31_120_2 = reservoir_state[120] <<< 2;
wire signed [31:0] shifted_state31_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state31_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state31_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state31_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state31_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state31_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state31_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state31_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state31_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state31_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state31_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state31_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state31_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state31_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state31_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state31_149_1 = reservoir_state[149] <<< 1;
wire signed [31:0] shifted_state31_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state31_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state31_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state31_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state31_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state31_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state31_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state31_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state31_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state31_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state31_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state31_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state31_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state31_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state31_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state31_179_2 = reservoir_state[179] <<< 2;
wire signed [31:0] shifted_state31_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state31_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state31_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state31_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state31_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state31_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state31_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state31_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state31_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state31_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state31_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state31_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state31_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state31_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state31_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state31_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state31_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state31_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state32_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state32_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state32_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state32_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state32_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state32_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state32_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state32_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state32_14_0 = reservoir_state[14] <<< 0;
wire signed [31:0] shifted_state32_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state32_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state32_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state32_39_0 = reservoir_state[39] <<< 0;
wire signed [31:0] shifted_state32_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state32_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state32_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state32_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state32_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state32_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state32_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state32_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state32_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state32_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state32_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state32_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state32_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state32_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state32_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state32_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state32_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state32_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state32_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state32_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state32_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state32_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state32_102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state32_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state32_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state32_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state32_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state32_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state32_124_3 = reservoir_state[124] <<< 3;
wire signed [31:0] shifted_state32_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state32_124_6 = reservoir_state[124] <<< 6;
wire signed [31:0] shifted_state32_124_7 = reservoir_state[124] <<< 7;
wire signed [31:0] shifted_state32_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state32_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state32_126_3 = reservoir_state[126] <<< 3;
wire signed [31:0] shifted_state32_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state32_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state32_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state32_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state32_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state32_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state32_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state32_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state32_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state32_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state32_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state32_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state32_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state32_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state32_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state32_161_0 = reservoir_state[161] <<< 0;
wire signed [31:0] shifted_state32_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state32_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state32_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state32_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state32_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state32_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state32_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state32_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state32_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state32_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state32_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state32_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state32_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state32_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state33_2_0 = reservoir_state[2] <<< 0;
wire signed [31:0] shifted_state33_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state33_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state33_2_3 = reservoir_state[2] <<< 3;
wire signed [31:0] shifted_state33_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state33_8_3 = reservoir_state[8] <<< 3;
wire signed [31:0] shifted_state33_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state33_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state33_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state33_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state33_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state33_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state33_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state33_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state33_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state33_17_4 = reservoir_state[17] <<< 4;
wire signed [31:0] shifted_state33_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state33_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state33_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state33_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state33_34_2 = reservoir_state[34] <<< 2;
wire signed [31:0] shifted_state33_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state33_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state33_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state33_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state33_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state33_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state33_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state33_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state33_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state33_51_6 = reservoir_state[51] <<< 6;
wire signed [31:0] shifted_state33_51_7 = reservoir_state[51] <<< 7;
wire signed [31:0] shifted_state33_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state33_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state33_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state33_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state33_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state33_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state33_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state33_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state33_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state33_79_5 = reservoir_state[79] <<< 5;
wire signed [31:0] shifted_state33_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state33_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state33_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state33_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state33_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state33_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state33_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state33_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state33_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state33_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state33_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state33_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state33_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state33_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state33_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state33_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state33_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state33_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state33_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state33_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state33_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state33_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state33_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state33_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state33_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state33_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state33_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state33_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state33_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state33_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state33_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state33_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state33_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state33_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state33_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state33_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state33_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state33_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state33_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state33_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state33_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state33_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state33_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state33_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state33_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state33_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state33_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state33_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state33_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state33_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state33_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state33_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state34_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state34_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state34_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state34_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state34_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state34_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state34_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state34_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state34_36_4 = reservoir_state[36] <<< 4;
wire signed [31:0] shifted_state34_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state34_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state34_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state34_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state34_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state34_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state34_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state34_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state34_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state34_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state34_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state34_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state34_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state34_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state34_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state34_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state34_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state34_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state34_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state34_90_1 = reservoir_state[90] <<< 1;
wire signed [31:0] shifted_state34_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state34_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state34_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state34_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state34_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state34_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state34_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state34_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state34_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state34_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state34_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state34_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state34_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state34_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state34_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state34_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state34_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state34_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state34_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state34_108_4 = reservoir_state[108] <<< 4;
wire signed [31:0] shifted_state34_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state34_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state34_120_2 = reservoir_state[120] <<< 2;
wire signed [31:0] shifted_state34_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state34_120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state34_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state34_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state34_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state34_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state34_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state34_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state34_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state34_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state34_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state34_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state34_148_6 = reservoir_state[148] <<< 6;
wire signed [31:0] shifted_state34_148_7 = reservoir_state[148] <<< 7;
wire signed [31:0] shifted_state34_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state34_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state34_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state34_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state34_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state34_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state34_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state34_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state34_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state34_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state34_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state34_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state34_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state34_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state34_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state34_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state34_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state34_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state35_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state35_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state35_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state35_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state35_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state35_23_5 = reservoir_state[23] <<< 5;
wire signed [31:0] shifted_state35_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state35_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state35_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state35_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state35_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state35_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state35_56_0 = reservoir_state[56] <<< 0;
wire signed [31:0] shifted_state35_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state35_56_5 = reservoir_state[56] <<< 5;
wire signed [31:0] shifted_state35_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state35_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state35_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state35_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state35_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state35_64_4 = reservoir_state[64] <<< 4;
wire signed [31:0] shifted_state35_64_6 = reservoir_state[64] <<< 6;
wire signed [31:0] shifted_state35_64_7 = reservoir_state[64] <<< 7;
wire signed [31:0] shifted_state35_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state35_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state35_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state35_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state35_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state35_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state35_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state35_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state35_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state35_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state35_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state35_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state35_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state35_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state35_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state35_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state35_102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state35_102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state35_102_7 = reservoir_state[102] <<< 7;
wire signed [31:0] shifted_state35_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state35_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state35_122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state35_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state35_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state35_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state35_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state35_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state35_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state35_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state35_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state35_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state35_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state35_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state35_145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state35_157_0 = reservoir_state[157] <<< 0;
wire signed [31:0] shifted_state35_157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state35_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state35_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state35_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state35_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state35_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state35_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state35_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state35_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state35_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state35_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state35_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state35_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state35_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state35_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state35_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state35_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state35_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state35_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state35_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state35_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state35_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state35_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state35_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state35_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state35_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state35_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state35_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state35_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state35_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state35_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state35_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state35_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state35_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state35_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state35_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state36_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state36_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state36_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state36_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state36_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state36_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state36_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state36_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state36_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state36_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state36_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state36_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state36_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state36_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state36_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state36_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state36_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state36_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state36_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state36_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state36_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state36_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state36_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state36_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state36_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state36_50_4 = reservoir_state[50] <<< 4;
wire signed [31:0] shifted_state36_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state36_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state36_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state36_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state36_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state36_70_4 = reservoir_state[70] <<< 4;
wire signed [31:0] shifted_state36_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state36_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state36_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state36_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state36_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state36_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state36_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state36_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state36_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state36_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state36_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state36_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state36_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state36_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state36_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state36_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state36_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state36_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state36_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state36_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state36_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state36_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state36_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state36_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state36_143_0 = reservoir_state[143] <<< 0;
wire signed [31:0] shifted_state36_143_3 = reservoir_state[143] <<< 3;
wire signed [31:0] shifted_state36_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state36_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state36_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state36_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state36_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state36_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state36_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state36_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state36_160_4 = reservoir_state[160] <<< 4;
wire signed [31:0] shifted_state36_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state36_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state36_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state36_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state36_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state36_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state36_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state36_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state36_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state36_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state36_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state36_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state37_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state37_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state37_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state37_33_4 = reservoir_state[33] <<< 4;
wire signed [31:0] shifted_state37_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state37_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state37_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state37_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state37_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state37_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state37_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state37_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state37_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state37_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state37_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state37_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state37_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state37_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state37_88_6 = reservoir_state[88] <<< 6;
wire signed [31:0] shifted_state37_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state37_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state37_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state37_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state37_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state37_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state37_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state37_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state37_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state37_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state37_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state37_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state37_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state37_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state37_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state37_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state37_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state37_158_0 = reservoir_state[158] <<< 0;
wire signed [31:0] shifted_state37_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state37_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state37_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state37_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state37_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state37_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state37_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state37_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state37_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state37_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state37_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state37_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state37_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state37_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state37_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state37_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state37_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state37_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state37_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state37_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state37_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state37_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state37_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state37_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state37_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state37_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state37_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state37_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state37_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state37_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state37_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state37_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state37_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state37_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state38_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state38_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state38_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state38_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state38_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state38_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state38_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state38_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state38_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state38_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state38_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state38_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state38_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state38_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state38_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state38_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state38_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state38_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state38_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state38_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state38_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state38_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state38_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state38_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state38_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state38_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state38_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state38_72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state38_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state38_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state38_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state38_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state38_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state38_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state38_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state38_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state38_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state38_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state38_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state38_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state38_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state38_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state38_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state38_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state38_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state38_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state38_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state38_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state38_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state38_103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state38_103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state38_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state38_120_2 = reservoir_state[120] <<< 2;
wire signed [31:0] shifted_state38_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state38_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state38_124_2 = reservoir_state[124] <<< 2;
wire signed [31:0] shifted_state38_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state38_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state38_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state38_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state38_135_3 = reservoir_state[135] <<< 3;
wire signed [31:0] shifted_state38_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state38_157_0 = reservoir_state[157] <<< 0;
wire signed [31:0] shifted_state38_157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state38_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state38_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state38_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state38_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state38_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state38_162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state38_162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state38_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state38_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state38_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state38_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state38_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state38_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state38_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state38_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state38_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state38_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state38_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state38_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state38_179_2 = reservoir_state[179] <<< 2;
wire signed [31:0] shifted_state38_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state39_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state39_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state39_1_3 = reservoir_state[1] <<< 3;
wire signed [31:0] shifted_state39_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state39_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state39_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state39_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state39_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state39_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state39_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state39_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state39_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state39_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state39_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state39_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state39_34_2 = reservoir_state[34] <<< 2;
wire signed [31:0] shifted_state39_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state39_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state39_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state39_69_1 = reservoir_state[69] <<< 1;
wire signed [31:0] shifted_state39_69_2 = reservoir_state[69] <<< 2;
wire signed [31:0] shifted_state39_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state39_69_5 = reservoir_state[69] <<< 5;
wire signed [31:0] shifted_state39_69_6 = reservoir_state[69] <<< 6;
wire signed [31:0] shifted_state39_69_7 = reservoir_state[69] <<< 7;
wire signed [31:0] shifted_state39_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state39_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state39_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state39_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state39_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state39_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state39_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state39_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state39_85_7 = reservoir_state[85] <<< 7;
wire signed [31:0] shifted_state39_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state39_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state39_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state39_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state39_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state39_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state39_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state39_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state39_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state39_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state39_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state39_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state39_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state39_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state39_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state39_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state39_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state39_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state39_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state39_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state39_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state39_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state39_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state39_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state39_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state39_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state39_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state39_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state39_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state39_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state39_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state39_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state39_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state39_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state39_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state39_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state39_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state39_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state39_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state39_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state39_161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state39_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state39_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state39_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state39_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state39_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state39_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state39_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state39_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state39_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state39_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state39_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state39_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state39_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state39_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state39_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state39_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state39_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state39_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state39_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state39_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state39_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state39_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state39_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state39_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state39_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state39_176_2 = reservoir_state[176] <<< 2;
wire signed [31:0] shifted_state39_176_4 = reservoir_state[176] <<< 4;
wire signed [31:0] shifted_state39_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state39_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state39_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state40_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state40_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state40_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state40_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state40_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state40_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state40_9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state40_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state40_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state40_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state40_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state40_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state40_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state40_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state40_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state40_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state40_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state40_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state40_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state40_23_5 = reservoir_state[23] <<< 5;
wire signed [31:0] shifted_state40_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state40_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state40_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state40_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state40_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state40_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state40_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state40_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state40_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state40_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state40_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state40_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state40_48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state40_48_5 = reservoir_state[48] <<< 5;
wire signed [31:0] shifted_state40_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state40_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state40_57_3 = reservoir_state[57] <<< 3;
wire signed [31:0] shifted_state40_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state40_75_3 = reservoir_state[75] <<< 3;
wire signed [31:0] shifted_state40_75_4 = reservoir_state[75] <<< 4;
wire signed [31:0] shifted_state40_75_5 = reservoir_state[75] <<< 5;
wire signed [31:0] shifted_state40_75_6 = reservoir_state[75] <<< 6;
wire signed [31:0] shifted_state40_75_7 = reservoir_state[75] <<< 7;
wire signed [31:0] shifted_state40_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state40_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state40_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state40_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state40_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state40_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state40_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state40_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state40_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state40_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state40_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state40_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state40_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state40_112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state40_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state40_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state40_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state40_119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state40_119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state40_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state40_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state40_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state40_120_5 = reservoir_state[120] <<< 5;
wire signed [31:0] shifted_state40_120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state40_120_7 = reservoir_state[120] <<< 7;
wire signed [31:0] shifted_state40_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state40_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state40_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state40_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state40_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state40_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state40_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state40_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state40_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state40_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state40_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state40_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state40_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state40_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state40_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state40_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state40_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state40_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state40_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state40_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state40_153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state40_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state40_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state40_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state40_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state40_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state40_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state40_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state40_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state40_156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state40_156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state40_156_6 = reservoir_state[156] <<< 6;
wire signed [31:0] shifted_state40_156_7 = reservoir_state[156] <<< 7;
wire signed [31:0] shifted_state40_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state40_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state40_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state40_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state41_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state41_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state41_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state41_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state41_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state41_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state41_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state41_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state41_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state41_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state41_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state41_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state41_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state41_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state41_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state41_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state41_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state41_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state41_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state41_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state41_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state41_53_3 = reservoir_state[53] <<< 3;
wire signed [31:0] shifted_state41_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state41_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state41_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state41_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state41_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state41_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state41_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state41_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state41_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state41_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state41_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state41_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state41_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state41_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state41_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state41_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state41_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state41_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state41_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state41_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state41_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state41_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state41_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state41_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state41_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state41_112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state41_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state41_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state41_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state41_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state41_147_5 = reservoir_state[147] <<< 5;
wire signed [31:0] shifted_state41_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state41_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state41_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state41_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state41_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state41_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state41_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state41_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state41_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state41_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state41_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state41_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state41_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state41_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state41_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state41_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state41_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state41_179_2 = reservoir_state[179] <<< 2;
wire signed [31:0] shifted_state41_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state41_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state41_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state41_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state41_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state41_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state41_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state41_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state41_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state42_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state42_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state42_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state42_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state42_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state42_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state42_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state42_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state42_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state42_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state42_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state42_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state42_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state42_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state42_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state42_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state42_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state42_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state42_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state42_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state42_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state42_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state42_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state42_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state42_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state42_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state42_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state42_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state42_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state42_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state42_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state42_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state42_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state42_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state42_143_0 = reservoir_state[143] <<< 0;
wire signed [31:0] shifted_state42_143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state42_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state42_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state42_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state42_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state42_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state42_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state42_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state42_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state42_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state42_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state42_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state42_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state43_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state43_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state43_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state43_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state43_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state43_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state43_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state43_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state43_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state43_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state43_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state43_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state43_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state43_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state43_93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state43_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state43_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state43_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state43_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state43_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state43_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state43_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state43_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state43_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state43_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state43_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state43_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state43_135_2 = reservoir_state[135] <<< 2;
wire signed [31:0] shifted_state43_135_4 = reservoir_state[135] <<< 4;
wire signed [31:0] shifted_state43_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state43_135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state43_135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state43_158_0 = reservoir_state[158] <<< 0;
wire signed [31:0] shifted_state43_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state43_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state43_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state43_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state43_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state43_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state43_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state43_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state43_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state43_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state44_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state44_3_1 = reservoir_state[3] <<< 1;
wire signed [31:0] shifted_state44_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state44_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state44_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state44_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state44_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state44_16_3 = reservoir_state[16] <<< 3;
wire signed [31:0] shifted_state44_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state44_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state44_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state44_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state44_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state44_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state44_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state44_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state44_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state44_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state44_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state44_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state44_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state44_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state44_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state44_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state44_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state44_68_1 = reservoir_state[68] <<< 1;
wire signed [31:0] shifted_state44_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state44_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state44_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state44_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state44_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state44_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state44_69_1 = reservoir_state[69] <<< 1;
wire signed [31:0] shifted_state44_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state44_69_5 = reservoir_state[69] <<< 5;
wire signed [31:0] shifted_state44_69_6 = reservoir_state[69] <<< 6;
wire signed [31:0] shifted_state44_69_7 = reservoir_state[69] <<< 7;
wire signed [31:0] shifted_state44_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state44_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state44_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state44_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state44_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state44_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state44_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state44_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state44_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state44_79_5 = reservoir_state[79] <<< 5;
wire signed [31:0] shifted_state44_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state44_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state44_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state44_87_2 = reservoir_state[87] <<< 2;
wire signed [31:0] shifted_state44_87_3 = reservoir_state[87] <<< 3;
wire signed [31:0] shifted_state44_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state44_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state44_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state44_91_1 = reservoir_state[91] <<< 1;
wire signed [31:0] shifted_state44_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state44_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state44_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state44_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state44_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state44_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state44_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state44_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state44_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state44_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state44_147_5 = reservoir_state[147] <<< 5;
wire signed [31:0] shifted_state44_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state44_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state44_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state44_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state44_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state44_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state44_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state44_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state44_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state44_186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state44_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state44_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state44_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state44_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state44_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state44_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state44_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state44_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state44_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state45_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state45_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state45_29_2 = reservoir_state[29] <<< 2;
wire signed [31:0] shifted_state45_29_3 = reservoir_state[29] <<< 3;
wire signed [31:0] shifted_state45_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state45_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state45_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state45_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state45_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state45_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state45_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state45_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state45_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state45_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state45_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state45_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state45_55_2 = reservoir_state[55] <<< 2;
wire signed [31:0] shifted_state45_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state45_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state45_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state45_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state45_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state45_58_2 = reservoir_state[58] <<< 2;
wire signed [31:0] shifted_state45_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state45_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state45_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state45_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state45_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state45_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state45_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state45_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state45_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state45_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state45_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state45_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state45_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state45_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state45_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state45_79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state45_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state45_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state45_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state45_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state45_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state45_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state45_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state45_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state45_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state45_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state45_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state45_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state45_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state45_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state45_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state45_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state45_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state45_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state45_91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state45_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state45_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state45_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state45_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state45_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state45_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state45_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state45_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state45_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state45_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state45_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state45_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state45_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state45_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state45_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state45_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state45_124_2 = reservoir_state[124] <<< 2;
wire signed [31:0] shifted_state45_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state45_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state45_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state45_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state45_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state45_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state45_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state45_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state45_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state45_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state45_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state45_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state45_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state45_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state45_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state45_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state45_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state45_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state45_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state45_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state45_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state45_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state45_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state45_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state45_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state45_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state45_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state45_197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state45_197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state45_197_5 = reservoir_state[197] <<< 5;
wire signed [31:0] shifted_state45_197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state45_197_7 = reservoir_state[197] <<< 7;
wire signed [31:0] shifted_state46_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state46_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state46_40_2 = reservoir_state[40] <<< 2;
wire signed [31:0] shifted_state46_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state46_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state46_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state46_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state46_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state46_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state46_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state46_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state46_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state46_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state46_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state46_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state46_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state46_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state46_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state46_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state46_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state46_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state46_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state46_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state46_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state46_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state46_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state46_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state46_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state46_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state46_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state46_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state46_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state46_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state46_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state46_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state46_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state46_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state46_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state46_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state46_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state46_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state46_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state46_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state46_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state46_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state46_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state46_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state46_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state46_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state46_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state46_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state46_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state46_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state46_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state46_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state46_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state46_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state46_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state46_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state46_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state46_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state46_146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state46_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state46_146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state46_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state46_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state46_147_1 = reservoir_state[147] <<< 1;
wire signed [31:0] shifted_state46_147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state46_147_6 = reservoir_state[147] <<< 6;
wire signed [31:0] shifted_state46_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state46_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state46_149_6 = reservoir_state[149] <<< 6;
wire signed [31:0] shifted_state46_149_7 = reservoir_state[149] <<< 7;
wire signed [31:0] shifted_state46_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state46_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state46_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state46_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state46_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state46_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state46_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state46_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state46_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state46_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state46_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state47_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state47_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state47_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state47_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state47_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state47_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state47_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state47_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state47_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state47_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state47_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state47_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state47_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state47_53_3 = reservoir_state[53] <<< 3;
wire signed [31:0] shifted_state47_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state47_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state47_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state47_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state47_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state47_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state47_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state47_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state47_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state47_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state47_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state47_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state47_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state47_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state47_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state47_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state47_73_1 = reservoir_state[73] <<< 1;
wire signed [31:0] shifted_state47_73_2 = reservoir_state[73] <<< 2;
wire signed [31:0] shifted_state47_73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state47_73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state47_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state47_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state47_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state47_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state47_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state47_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state47_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state47_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state47_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state47_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state47_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state47_98_5 = reservoir_state[98] <<< 5;
wire signed [31:0] shifted_state47_98_6 = reservoir_state[98] <<< 6;
wire signed [31:0] shifted_state47_98_7 = reservoir_state[98] <<< 7;
wire signed [31:0] shifted_state47_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state47_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state47_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state47_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state47_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state47_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state47_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state47_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state47_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state47_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state47_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state47_146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state47_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state47_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state47_146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state47_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state47_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state47_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state47_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state47_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state47_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state47_159_0 = reservoir_state[159] <<< 0;
wire signed [31:0] shifted_state47_159_5 = reservoir_state[159] <<< 5;
wire signed [31:0] shifted_state47_185_2 = reservoir_state[185] <<< 2;
wire signed [31:0] shifted_state47_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state47_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state47_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state47_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state47_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state47_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state47_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state47_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state47_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state48_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state48_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state48_8_5 = reservoir_state[8] <<< 5;
wire signed [31:0] shifted_state48_8_6 = reservoir_state[8] <<< 6;
wire signed [31:0] shifted_state48_8_7 = reservoir_state[8] <<< 7;
wire signed [31:0] shifted_state48_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state48_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state48_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state48_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state48_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state48_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state48_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state48_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state48_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state48_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state48_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state48_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state48_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state48_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state48_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state48_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state48_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state48_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state48_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state48_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state48_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state48_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state48_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state48_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state48_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state48_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state48_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state48_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state48_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state48_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state48_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state48_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state48_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state48_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state48_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state48_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state48_94_2 = reservoir_state[94] <<< 2;
wire signed [31:0] shifted_state48_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state48_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state48_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state48_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state48_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state48_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state48_102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state48_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state48_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state48_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state48_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state48_125_2 = reservoir_state[125] <<< 2;
wire signed [31:0] shifted_state48_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state48_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state48_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state48_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state48_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state48_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state48_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state48_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state48_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state48_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state48_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state48_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state48_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state48_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state48_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state48_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state48_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state48_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state48_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state48_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state48_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state48_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state48_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state48_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state48_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state48_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state48_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state48_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state48_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state48_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state48_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state48_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state48_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state48_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state48_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state48_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state48_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state48_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state48_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state48_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state48_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state48_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state48_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state48_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state48_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state48_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state48_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state49_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state49_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state49_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state49_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state49_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state49_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state49_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state49_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state49_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state49_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state49_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state49_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state49_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state49_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state49_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state49_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state49_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state49_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state49_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state49_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state49_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state49_74_3 = reservoir_state[74] <<< 3;
wire signed [31:0] shifted_state49_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state49_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state49_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state49_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state49_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state49_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state49_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state49_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state49_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state49_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state49_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state49_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state49_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state49_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state49_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state49_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state49_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state49_157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state49_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state49_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state49_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state49_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state49_159_0 = reservoir_state[159] <<< 0;
wire signed [31:0] shifted_state49_159_1 = reservoir_state[159] <<< 1;
wire signed [31:0] shifted_state49_159_2 = reservoir_state[159] <<< 2;
wire signed [31:0] shifted_state50_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state50_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state50_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state50_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state50_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state50_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state50_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state50_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state50_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state50_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state50_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state50_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state50_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state50_66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state50_66_2 = reservoir_state[66] <<< 2;
wire signed [31:0] shifted_state50_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state50_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state50_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state50_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state50_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state50_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state50_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state50_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state50_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state50_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state50_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state50_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state50_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state50_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state50_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state50_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state50_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state50_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state50_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state50_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state50_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state50_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state50_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state50_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state50_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state50_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state50_110_1 = reservoir_state[110] <<< 1;
wire signed [31:0] shifted_state50_110_2 = reservoir_state[110] <<< 2;
wire signed [31:0] shifted_state50_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state50_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state50_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state50_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state50_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state50_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state50_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state50_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state50_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state50_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state50_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state50_161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state50_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state50_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state50_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state50_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state50_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state50_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state50_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state50_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state50_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state50_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state50_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state50_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state50_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state50_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state50_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state50_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state50_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state50_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state50_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state50_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state50_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state51_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state51_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state51_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state51_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state51_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state51_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state51_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state51_58_2 = reservoir_state[58] <<< 2;
wire signed [31:0] shifted_state51_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state51_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state51_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state51_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state51_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state51_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state51_66_2 = reservoir_state[66] <<< 2;
wire signed [31:0] shifted_state51_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state51_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state51_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state51_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state51_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state51_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state51_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state51_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state51_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state51_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state51_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state51_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state51_108_4 = reservoir_state[108] <<< 4;
wire signed [31:0] shifted_state51_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state51_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state51_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state51_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state51_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state51_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state51_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state51_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state51_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state51_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state51_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state51_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state51_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state51_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state51_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state51_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state51_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state51_199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state52_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state52_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state52_9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state52_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state52_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state52_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state52_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state52_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state52_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state52_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state52_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state52_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state52_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state52_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state52_48_5 = reservoir_state[48] <<< 5;
wire signed [31:0] shifted_state52_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state52_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state52_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state52_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state52_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state52_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state52_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state52_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state52_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state52_79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state52_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state52_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state52_79_5 = reservoir_state[79] <<< 5;
wire signed [31:0] shifted_state52_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state52_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state52_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state52_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state52_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state52_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state52_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state52_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state52_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state52_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state52_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state52_112_3 = reservoir_state[112] <<< 3;
wire signed [31:0] shifted_state52_119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state52_119_2 = reservoir_state[119] <<< 2;
wire signed [31:0] shifted_state52_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state52_119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state52_119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state52_142_0 = reservoir_state[142] <<< 0;
wire signed [31:0] shifted_state52_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state52_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state52_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state52_144_0 = reservoir_state[144] <<< 0;
wire signed [31:0] shifted_state52_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state52_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state52_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state52_151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state52_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state52_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state52_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state52_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state52_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state52_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state52_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state52_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state52_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state52_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state52_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state52_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state52_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state52_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state52_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state52_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state52_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state52_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state52_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state52_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state52_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state53_1_3 = reservoir_state[1] <<< 3;
wire signed [31:0] shifted_state53_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state53_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state53_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state53_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state53_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state53_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state53_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state53_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state53_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state53_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state53_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state53_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state53_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state53_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state53_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state53_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state53_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state53_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state53_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state53_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state53_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state53_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state53_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state53_27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state53_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state53_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state53_27_4 = reservoir_state[27] <<< 4;
wire signed [31:0] shifted_state53_27_5 = reservoir_state[27] <<< 5;
wire signed [31:0] shifted_state53_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state53_29_2 = reservoir_state[29] <<< 2;
wire signed [31:0] shifted_state53_29_3 = reservoir_state[29] <<< 3;
wire signed [31:0] shifted_state53_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state53_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state53_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state53_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state53_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state53_30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state53_30_4 = reservoir_state[30] <<< 4;
wire signed [31:0] shifted_state53_30_5 = reservoir_state[30] <<< 5;
wire signed [31:0] shifted_state53_30_6 = reservoir_state[30] <<< 6;
wire signed [31:0] shifted_state53_30_7 = reservoir_state[30] <<< 7;
wire signed [31:0] shifted_state53_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state53_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state53_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state53_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state53_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state53_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state53_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state53_64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state53_64_6 = reservoir_state[64] <<< 6;
wire signed [31:0] shifted_state53_64_7 = reservoir_state[64] <<< 7;
wire signed [31:0] shifted_state53_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state53_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state53_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state53_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state53_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state53_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state53_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state53_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state53_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state53_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state53_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state53_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state53_142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state53_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state53_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state53_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state53_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state53_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state53_148_6 = reservoir_state[148] <<< 6;
wire signed [31:0] shifted_state53_148_7 = reservoir_state[148] <<< 7;
wire signed [31:0] shifted_state53_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state53_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state53_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state53_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state53_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state53_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state53_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state53_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state53_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state53_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state53_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state53_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state53_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state53_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state53_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state53_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state53_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state53_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state53_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state53_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state54_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state54_23_4 = reservoir_state[23] <<< 4;
wire signed [31:0] shifted_state54_23_5 = reservoir_state[23] <<< 5;
wire signed [31:0] shifted_state54_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state54_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state54_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state54_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state54_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state54_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state54_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state54_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state54_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state54_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state54_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state54_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state54_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state54_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state54_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state54_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state54_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state54_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state54_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state54_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state54_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state54_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state54_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state54_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state54_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state54_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state54_70_2 = reservoir_state[70] <<< 2;
wire signed [31:0] shifted_state54_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state54_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state54_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state54_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state54_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state54_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state54_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state54_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state54_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state54_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state54_110_1 = reservoir_state[110] <<< 1;
wire signed [31:0] shifted_state54_110_4 = reservoir_state[110] <<< 4;
wire signed [31:0] shifted_state54_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state54_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state54_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state54_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state54_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state54_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state54_115_3 = reservoir_state[115] <<< 3;
wire signed [31:0] shifted_state54_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state54_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state54_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state54_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state54_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state54_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state54_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state54_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state54_156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state54_156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state54_156_6 = reservoir_state[156] <<< 6;
wire signed [31:0] shifted_state54_156_7 = reservoir_state[156] <<< 7;
wire signed [31:0] shifted_state54_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state54_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state54_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state54_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state54_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state54_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state54_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state54_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state54_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state54_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state54_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state54_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state54_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state54_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state54_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state54_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state54_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state54_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state54_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state54_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state55_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state55_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state55_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state55_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state55_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state55_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state55_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state55_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state55_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state55_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state55_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state55_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state55_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state55_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state55_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state55_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state55_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state55_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state55_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state55_125_2 = reservoir_state[125] <<< 2;
wire signed [31:0] shifted_state55_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state55_125_5 = reservoir_state[125] <<< 5;
wire signed [31:0] shifted_state55_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state55_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state55_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state55_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state55_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state55_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state55_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state55_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state55_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state55_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state55_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state55_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state55_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state55_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state55_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state55_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state55_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state55_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state55_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state55_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state55_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state55_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state55_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state55_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state55_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state55_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state55_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state55_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state55_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state55_169_2 = reservoir_state[169] <<< 2;
wire signed [31:0] shifted_state55_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state55_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state55_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state55_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state55_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state55_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state55_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state55_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state55_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state55_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state55_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state55_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state55_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state55_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state56_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state56_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state56_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state56_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state56_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state56_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state56_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state56_12_0 = reservoir_state[12] <<< 0;
wire signed [31:0] shifted_state56_12_5 = reservoir_state[12] <<< 5;
wire signed [31:0] shifted_state56_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state56_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state56_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state56_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state56_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state56_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state56_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state56_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state56_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state56_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state56_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state56_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state56_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state56_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state56_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state56_66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state56_66_2 = reservoir_state[66] <<< 2;
wire signed [31:0] shifted_state56_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state56_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state56_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state56_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state56_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state56_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state56_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state56_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state56_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state56_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state56_90_0 = reservoir_state[90] <<< 0;
wire signed [31:0] shifted_state56_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state56_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state56_90_4 = reservoir_state[90] <<< 4;
wire signed [31:0] shifted_state56_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state56_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state56_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state56_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state56_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state56_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state56_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state56_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state56_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state56_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state56_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state56_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state56_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state56_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state56_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state56_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state56_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state56_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state56_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state56_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state56_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state56_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state56_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state56_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state56_120_2 = reservoir_state[120] <<< 2;
wire signed [31:0] shifted_state56_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state56_120_5 = reservoir_state[120] <<< 5;
wire signed [31:0] shifted_state56_120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state56_120_7 = reservoir_state[120] <<< 7;
wire signed [31:0] shifted_state56_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state56_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state56_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state56_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state56_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state56_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state56_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state56_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state56_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state56_157_0 = reservoir_state[157] <<< 0;
wire signed [31:0] shifted_state56_157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state56_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state56_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state56_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state56_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state56_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state56_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state56_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state57_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state57_34_2 = reservoir_state[34] <<< 2;
wire signed [31:0] shifted_state57_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state57_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state57_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state57_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state57_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state57_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state57_55_2 = reservoir_state[55] <<< 2;
wire signed [31:0] shifted_state57_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state57_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state57_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state57_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state57_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state57_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state57_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state57_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state57_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state57_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state57_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state57_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state57_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state57_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state57_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state57_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state57_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state57_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state57_115_3 = reservoir_state[115] <<< 3;
wire signed [31:0] shifted_state57_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state57_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state57_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state57_142_0 = reservoir_state[142] <<< 0;
wire signed [31:0] shifted_state57_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state57_142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state57_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state57_147_1 = reservoir_state[147] <<< 1;
wire signed [31:0] shifted_state57_147_3 = reservoir_state[147] <<< 3;
wire signed [31:0] shifted_state57_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state57_154_0 = reservoir_state[154] <<< 0;
wire signed [31:0] shifted_state57_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state57_154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state57_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state57_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state57_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state57_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state57_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state57_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state57_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state57_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state57_156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state57_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state57_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state57_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state57_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state57_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state57_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state57_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state57_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state57_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state57_167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state57_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state57_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state57_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state57_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state57_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state57_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state57_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state57_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state57_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state57_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state57_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state57_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state57_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state58_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state58_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state58_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state58_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state58_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state58_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state58_29_3 = reservoir_state[29] <<< 3;
wire signed [31:0] shifted_state58_29_5 = reservoir_state[29] <<< 5;
wire signed [31:0] shifted_state58_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state58_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state58_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state58_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state58_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state58_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state58_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state58_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state58_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state58_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state58_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state58_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state58_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state58_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state58_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state58_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state58_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state58_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state58_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state58_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state58_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state58_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state58_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state58_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state58_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state58_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state58_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state58_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state58_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state58_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state58_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state58_98_6 = reservoir_state[98] <<< 6;
wire signed [31:0] shifted_state58_98_7 = reservoir_state[98] <<< 7;
wire signed [31:0] shifted_state58_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state58_110_0 = reservoir_state[110] <<< 0;
wire signed [31:0] shifted_state58_110_1 = reservoir_state[110] <<< 1;
wire signed [31:0] shifted_state58_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state58_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state58_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state58_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state58_137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state58_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state58_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state58_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state58_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state58_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state58_160_4 = reservoir_state[160] <<< 4;
wire signed [31:0] shifted_state58_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state58_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state58_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state58_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state58_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state58_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state58_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state58_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state58_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state59_15_0 = reservoir_state[15] <<< 0;
wire signed [31:0] shifted_state59_15_1 = reservoir_state[15] <<< 1;
wire signed [31:0] shifted_state59_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state59_15_3 = reservoir_state[15] <<< 3;
wire signed [31:0] shifted_state59_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state59_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state59_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state59_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state59_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state59_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state59_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state59_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state59_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state59_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state59_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state59_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state59_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state59_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state59_90_4 = reservoir_state[90] <<< 4;
wire signed [31:0] shifted_state59_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state59_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state59_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state59_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state59_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state59_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state59_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state59_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state59_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state59_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state59_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state59_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state59_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state59_115_4 = reservoir_state[115] <<< 4;
wire signed [31:0] shifted_state59_115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state59_115_6 = reservoir_state[115] <<< 6;
wire signed [31:0] shifted_state59_115_7 = reservoir_state[115] <<< 7;
wire signed [31:0] shifted_state59_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state59_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state59_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state59_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state59_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state59_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state59_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state59_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state59_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state59_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state59_136_2 = reservoir_state[136] <<< 2;
wire signed [31:0] shifted_state59_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state59_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state59_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state59_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state59_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state59_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state59_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state59_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state59_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state59_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state59_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state59_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state59_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state59_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state59_194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state59_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state59_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state59_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state59_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state59_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state59_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state59_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state59_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state60_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state60_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state60_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state60_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state60_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state60_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state60_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state60_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state60_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state60_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state60_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state60_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state60_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state60_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state60_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state60_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state60_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state60_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state60_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state60_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state60_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state60_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state60_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state60_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state60_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state60_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state60_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state60_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state60_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state60_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state60_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state60_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state60_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state60_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state60_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state60_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state60_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state60_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state60_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state60_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state60_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state60_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state60_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state60_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state60_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state60_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state60_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state60_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state60_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state60_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state60_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state60_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state60_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state60_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state60_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state60_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state60_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state60_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state60_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state60_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state60_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state60_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state60_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state60_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state60_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state60_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state60_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state60_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state60_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state60_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state60_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state60_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state60_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state60_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state60_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state60_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state60_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state60_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state60_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state60_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state60_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state60_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state60_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state61_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state61_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state61_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state61_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state61_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state61_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state61_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state61_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state61_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state61_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state61_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state61_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state61_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state61_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state61_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state61_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state61_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state61_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state61_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state61_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state61_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state61_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state61_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state61_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state61_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state61_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state61_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state61_84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state61_84_5 = reservoir_state[84] <<< 5;
wire signed [31:0] shifted_state61_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state61_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state61_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state61_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state61_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state61_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state61_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state61_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state61_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state61_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state61_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state61_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state61_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state61_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state61_117_5 = reservoir_state[117] <<< 5;
wire signed [31:0] shifted_state61_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state61_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state61_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state61_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state61_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state61_119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state61_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state61_119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state61_119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state61_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state61_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state61_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state61_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state61_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state61_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state61_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state61_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state61_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state61_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state61_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state61_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state61_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state61_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state61_142_0 = reservoir_state[142] <<< 0;
wire signed [31:0] shifted_state61_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state61_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state61_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state61_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state61_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state61_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state61_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state61_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state61_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state61_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state61_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state61_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state61_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state61_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state61_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state61_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state61_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state61_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state61_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state61_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state61_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state62_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state62_9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state62_14_0 = reservoir_state[14] <<< 0;
wire signed [31:0] shifted_state62_14_3 = reservoir_state[14] <<< 3;
wire signed [31:0] shifted_state62_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state62_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state62_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state62_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state62_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state62_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state62_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state62_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state62_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state62_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state62_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state62_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state62_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state62_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state62_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state62_47_5 = reservoir_state[47] <<< 5;
wire signed [31:0] shifted_state62_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state62_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state62_67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state62_67_1 = reservoir_state[67] <<< 1;
wire signed [31:0] shifted_state62_67_2 = reservoir_state[67] <<< 2;
wire signed [31:0] shifted_state62_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state62_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state62_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state62_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state62_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state62_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state62_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state62_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state62_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state62_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state62_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state62_134_0 = reservoir_state[134] <<< 0;
wire signed [31:0] shifted_state62_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state62_134_5 = reservoir_state[134] <<< 5;
wire signed [31:0] shifted_state62_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state62_134_7 = reservoir_state[134] <<< 7;
wire signed [31:0] shifted_state62_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state62_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state62_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state62_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state62_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state62_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state62_143_0 = reservoir_state[143] <<< 0;
wire signed [31:0] shifted_state62_143_2 = reservoir_state[143] <<< 2;
wire signed [31:0] shifted_state62_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state62_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state62_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state62_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state62_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state62_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state62_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state62_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state62_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state62_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state62_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state62_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state62_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state62_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state62_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state62_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state62_189_6 = reservoir_state[189] <<< 6;
wire signed [31:0] shifted_state62_189_7 = reservoir_state[189] <<< 7;
wire signed [31:0] shifted_state63_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state63_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state63_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state63_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state63_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state63_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state63_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state63_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state63_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state63_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state63_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state63_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state63_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state63_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state63_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state63_43_1 = reservoir_state[43] <<< 1;
wire signed [31:0] shifted_state63_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state63_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state63_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state63_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state63_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state63_73_5 = reservoir_state[73] <<< 5;
wire signed [31:0] shifted_state63_73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state63_73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state63_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state63_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state63_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state63_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state63_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state63_91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state63_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state63_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state63_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state63_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state63_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state63_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state63_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state63_92_6 = reservoir_state[92] <<< 6;
wire signed [31:0] shifted_state63_92_7 = reservoir_state[92] <<< 7;
wire signed [31:0] shifted_state63_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state63_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state63_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state63_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state63_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state63_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state63_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state63_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state63_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state63_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state63_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state63_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state63_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state63_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state63_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state63_128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state63_128_2 = reservoir_state[128] <<< 2;
wire signed [31:0] shifted_state63_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state63_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state63_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state63_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state63_131_2 = reservoir_state[131] <<< 2;
wire signed [31:0] shifted_state63_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state63_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state63_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state63_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state63_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state63_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state63_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state63_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state63_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state63_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state63_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state63_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state63_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state63_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state63_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state63_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state63_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state63_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state63_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state63_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state63_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state63_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state63_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state63_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state63_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state64_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state64_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state64_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state64_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state64_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state64_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state64_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state64_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state64_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state64_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state64_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state64_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state64_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state64_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state64_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state64_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state64_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state64_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state64_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state64_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state64_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state64_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state64_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state64_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state64_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state64_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state64_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state64_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state64_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state64_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state64_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state64_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state64_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state64_98_6 = reservoir_state[98] <<< 6;
wire signed [31:0] shifted_state64_98_7 = reservoir_state[98] <<< 7;
wire signed [31:0] shifted_state64_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state64_103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state64_103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state64_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state64_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state64_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state64_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state64_122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state64_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state64_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state64_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state64_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state64_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state64_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state64_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state64_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state64_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state64_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state64_128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state64_128_3 = reservoir_state[128] <<< 3;
wire signed [31:0] shifted_state64_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state64_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state64_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state64_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state64_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state64_134_0 = reservoir_state[134] <<< 0;
wire signed [31:0] shifted_state64_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state64_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state64_134_4 = reservoir_state[134] <<< 4;
wire signed [31:0] shifted_state64_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state64_134_7 = reservoir_state[134] <<< 7;
wire signed [31:0] shifted_state64_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state64_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state64_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state64_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state64_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state64_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state64_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state64_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state64_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state64_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state64_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state64_181_3 = reservoir_state[181] <<< 3;
wire signed [31:0] shifted_state64_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state64_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state64_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state64_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state64_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state64_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state64_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state64_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state64_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state64_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state65_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state65_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state65_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state65_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state65_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state65_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state65_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state65_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state65_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state65_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state65_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state65_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state65_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state65_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state65_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state65_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state65_13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state65_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state65_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state65_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state65_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state65_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state65_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state65_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state65_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state65_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state65_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state65_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state65_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state65_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state65_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state65_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state65_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state65_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state65_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state65_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state65_110_0 = reservoir_state[110] <<< 0;
wire signed [31:0] shifted_state65_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state65_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state65_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state65_111_4 = reservoir_state[111] <<< 4;
wire signed [31:0] shifted_state65_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state65_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state65_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state65_119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state65_119_2 = reservoir_state[119] <<< 2;
wire signed [31:0] shifted_state65_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state65_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state65_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state65_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state65_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state65_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state65_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state65_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state65_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state65_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state65_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state65_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state65_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state65_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state65_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state65_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state65_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state65_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state65_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state65_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state65_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state65_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state65_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state66_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state66_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state66_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state66_15_0 = reservoir_state[15] <<< 0;
wire signed [31:0] shifted_state66_15_1 = reservoir_state[15] <<< 1;
wire signed [31:0] shifted_state66_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state66_15_4 = reservoir_state[15] <<< 4;
wire signed [31:0] shifted_state66_15_6 = reservoir_state[15] <<< 6;
wire signed [31:0] shifted_state66_15_7 = reservoir_state[15] <<< 7;
wire signed [31:0] shifted_state66_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state66_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state66_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state66_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state66_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state66_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state66_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state66_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state66_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state66_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state66_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state66_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state66_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state66_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state66_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state66_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state66_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state66_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state66_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state66_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state66_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state66_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state66_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state66_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state66_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state66_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state66_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state66_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state66_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state66_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state66_115_4 = reservoir_state[115] <<< 4;
wire signed [31:0] shifted_state66_117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state66_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state66_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state66_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state66_119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state66_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state66_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state66_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state66_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state66_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state66_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state66_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state66_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state66_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state66_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state66_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state66_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state66_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state66_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state66_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state66_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state66_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state67_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state67_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state67_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state67_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state67_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state67_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state67_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state67_5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state67_5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state67_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state67_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state67_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state67_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state67_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state67_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state67_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state67_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state67_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state67_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state67_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state67_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state67_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state67_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state67_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state67_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state67_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state67_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state67_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state67_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state67_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state67_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state67_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state67_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state67_64_4 = reservoir_state[64] <<< 4;
wire signed [31:0] shifted_state67_64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state67_64_6 = reservoir_state[64] <<< 6;
wire signed [31:0] shifted_state67_64_7 = reservoir_state[64] <<< 7;
wire signed [31:0] shifted_state67_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state67_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state67_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state67_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state67_90_0 = reservoir_state[90] <<< 0;
wire signed [31:0] shifted_state67_90_1 = reservoir_state[90] <<< 1;
wire signed [31:0] shifted_state67_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state67_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state67_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state67_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state67_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state67_120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state67_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state67_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state67_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state67_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state67_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state67_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state67_144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state67_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state67_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state67_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state67_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state67_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state67_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state67_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state67_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state67_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state67_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state67_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state67_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state67_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state67_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state67_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state67_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state67_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state67_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state68_8_1 = reservoir_state[8] <<< 1;
wire signed [31:0] shifted_state68_8_3 = reservoir_state[8] <<< 3;
wire signed [31:0] shifted_state68_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state68_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state68_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state68_23_5 = reservoir_state[23] <<< 5;
wire signed [31:0] shifted_state68_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state68_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state68_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state68_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state68_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state68_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state68_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state68_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state68_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state68_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state68_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state68_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state68_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state68_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state68_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state68_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state68_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state68_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state68_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state68_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state68_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state68_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state68_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state68_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state68_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state68_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state68_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state68_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state68_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state68_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state68_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state68_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state68_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state68_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state68_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state68_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state68_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state68_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state68_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state68_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state68_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state68_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state68_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state68_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state68_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state68_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state68_148_6 = reservoir_state[148] <<< 6;
wire signed [31:0] shifted_state68_148_7 = reservoir_state[148] <<< 7;
wire signed [31:0] shifted_state68_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state68_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state68_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state68_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state68_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state68_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state68_159_2 = reservoir_state[159] <<< 2;
wire signed [31:0] shifted_state68_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state68_159_4 = reservoir_state[159] <<< 4;
wire signed [31:0] shifted_state68_159_6 = reservoir_state[159] <<< 6;
wire signed [31:0] shifted_state68_159_7 = reservoir_state[159] <<< 7;
wire signed [31:0] shifted_state68_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state68_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state68_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state68_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state68_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state68_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state68_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state69_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state69_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state69_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state69_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state69_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state69_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state69_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state69_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state69_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state69_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state69_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state69_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state69_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state69_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state69_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state69_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state69_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state69_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state69_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state69_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state69_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state69_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state69_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state69_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state69_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state69_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state69_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state69_49_3 = reservoir_state[49] <<< 3;
wire signed [31:0] shifted_state69_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state69_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state69_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state69_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state69_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state69_64_4 = reservoir_state[64] <<< 4;
wire signed [31:0] shifted_state69_64_6 = reservoir_state[64] <<< 6;
wire signed [31:0] shifted_state69_64_7 = reservoir_state[64] <<< 7;
wire signed [31:0] shifted_state69_74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state69_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state69_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state69_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state69_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state69_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state69_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state69_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state69_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state69_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state69_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state69_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state69_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state69_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state69_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state69_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state69_111_4 = reservoir_state[111] <<< 4;
wire signed [31:0] shifted_state69_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state69_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state69_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state69_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state69_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state69_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state69_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state69_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state69_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state69_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state69_148_6 = reservoir_state[148] <<< 6;
wire signed [31:0] shifted_state69_148_7 = reservoir_state[148] <<< 7;
wire signed [31:0] shifted_state69_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state69_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state69_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state69_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state69_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state69_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state69_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state69_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state69_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state70_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state70_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state70_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state70_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state70_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state70_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state70_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state70_66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state70_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state70_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state70_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state70_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state70_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state70_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state70_118_3 = reservoir_state[118] <<< 3;
wire signed [31:0] shifted_state70_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state70_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state70_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state70_126_3 = reservoir_state[126] <<< 3;
wire signed [31:0] shifted_state70_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state70_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state70_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state70_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state70_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state70_128_2 = reservoir_state[128] <<< 2;
wire signed [31:0] shifted_state70_128_5 = reservoir_state[128] <<< 5;
wire signed [31:0] shifted_state70_128_6 = reservoir_state[128] <<< 6;
wire signed [31:0] shifted_state70_128_7 = reservoir_state[128] <<< 7;
wire signed [31:0] shifted_state70_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state70_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state70_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state70_162_0 = reservoir_state[162] <<< 0;
wire signed [31:0] shifted_state70_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state70_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state70_162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state70_162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state70_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state70_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state70_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state70_182_1 = reservoir_state[182] <<< 1;
wire signed [31:0] shifted_state70_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state70_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state70_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state70_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state70_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state70_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state70_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state70_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state70_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state70_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state70_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state70_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state70_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state71_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state71_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state71_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state71_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state71_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state71_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state71_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state71_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state71_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state71_47_4 = reservoir_state[47] <<< 4;
wire signed [31:0] shifted_state71_47_5 = reservoir_state[47] <<< 5;
wire signed [31:0] shifted_state71_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state71_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state71_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state71_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state71_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state71_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state71_90_0 = reservoir_state[90] <<< 0;
wire signed [31:0] shifted_state71_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state71_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state71_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state71_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state71_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state71_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state71_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state71_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state71_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state71_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state71_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state71_103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state71_103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state71_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state71_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state71_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state71_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state71_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state71_151_4 = reservoir_state[151] <<< 4;
wire signed [31:0] shifted_state71_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state71_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state71_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state71_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state71_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state71_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state71_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state71_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state71_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state71_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state71_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state71_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state71_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state71_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state71_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state71_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state71_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state71_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state71_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state72_2_0 = reservoir_state[2] <<< 0;
wire signed [31:0] shifted_state72_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state72_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state72_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state72_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state72_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state72_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state72_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state72_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state72_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state72_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state72_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state72_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state72_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state72_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state72_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state72_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state72_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state72_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state72_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state72_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state72_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state72_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state72_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state72_66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state72_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state72_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state72_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state72_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state72_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state72_69_1 = reservoir_state[69] <<< 1;
wire signed [31:0] shifted_state72_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state72_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state72_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state72_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state72_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state72_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state72_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state72_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state72_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state72_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state72_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state72_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state72_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state72_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state72_102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state72_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state72_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state72_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state72_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state72_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state72_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state72_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state72_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state72_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state72_125_4 = reservoir_state[125] <<< 4;
wire signed [31:0] shifted_state72_125_5 = reservoir_state[125] <<< 5;
wire signed [31:0] shifted_state72_125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state72_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state72_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state72_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state72_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state72_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state72_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state72_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state72_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state72_143_0 = reservoir_state[143] <<< 0;
wire signed [31:0] shifted_state72_143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state72_143_3 = reservoir_state[143] <<< 3;
wire signed [31:0] shifted_state72_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state72_143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state72_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state72_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state72_144_0 = reservoir_state[144] <<< 0;
wire signed [31:0] shifted_state72_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state72_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state72_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state72_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state72_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state72_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state72_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state72_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state72_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state72_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state72_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state72_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state72_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state72_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state72_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state72_186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state72_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state73_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state73_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state73_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state73_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state73_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state73_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state73_43_1 = reservoir_state[43] <<< 1;
wire signed [31:0] shifted_state73_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state73_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state73_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state73_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state73_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state73_52_0 = reservoir_state[52] <<< 0;
wire signed [31:0] shifted_state73_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state73_70_2 = reservoir_state[70] <<< 2;
wire signed [31:0] shifted_state73_70_4 = reservoir_state[70] <<< 4;
wire signed [31:0] shifted_state73_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state73_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state73_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state73_72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state73_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state73_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state73_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state73_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state73_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state73_110_0 = reservoir_state[110] <<< 0;
wire signed [31:0] shifted_state73_110_2 = reservoir_state[110] <<< 2;
wire signed [31:0] shifted_state73_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state73_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state73_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state73_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state73_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state73_114_1 = reservoir_state[114] <<< 1;
wire signed [31:0] shifted_state73_114_2 = reservoir_state[114] <<< 2;
wire signed [31:0] shifted_state73_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state73_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state73_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state73_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state73_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state73_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state73_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state73_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state73_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state73_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state73_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state73_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state73_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state73_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state73_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state73_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state73_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state73_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state73_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state73_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state73_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state73_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state73_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state73_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state73_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state73_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state73_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state73_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state73_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state73_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state73_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state73_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state73_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state73_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state73_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state73_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state73_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state73_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state73_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state73_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state73_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state73_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state73_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state73_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state73_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state73_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state73_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state73_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state73_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state73_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state73_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state73_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state73_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state73_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state74_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state74_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state74_6_3 = reservoir_state[6] <<< 3;
wire signed [31:0] shifted_state74_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state74_13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state74_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state74_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state74_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state74_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state74_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state74_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state74_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state74_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state74_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state74_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state74_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state74_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state74_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state74_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state74_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state74_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state74_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state74_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state74_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state74_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state74_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state74_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state74_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state74_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state74_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state74_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state74_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state74_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state74_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state74_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state74_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state74_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state74_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state74_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state74_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state74_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state74_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state74_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state74_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state74_85_7 = reservoir_state[85] <<< 7;
wire signed [31:0] shifted_state74_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state74_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state74_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state74_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state74_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state74_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state74_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state74_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state74_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state74_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state74_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state74_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state74_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state74_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state74_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state74_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state74_98_5 = reservoir_state[98] <<< 5;
wire signed [31:0] shifted_state74_98_7 = reservoir_state[98] <<< 7;
wire signed [31:0] shifted_state74_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state74_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state74_118_3 = reservoir_state[118] <<< 3;
wire signed [31:0] shifted_state74_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state74_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state74_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state74_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state74_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state74_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state74_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state74_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state74_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state74_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state74_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state74_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state74_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state74_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state74_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state74_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state74_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state74_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state74_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state74_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state74_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state74_149_2 = reservoir_state[149] <<< 2;
wire signed [31:0] shifted_state74_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state74_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state74_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state74_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state74_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state74_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state74_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state74_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state74_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state74_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state74_176_0 = reservoir_state[176] <<< 0;
wire signed [31:0] shifted_state74_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state74_176_3 = reservoir_state[176] <<< 3;
wire signed [31:0] shifted_state74_176_5 = reservoir_state[176] <<< 5;
wire signed [31:0] shifted_state74_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state74_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state74_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state74_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state74_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state74_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state75_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state75_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state75_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state75_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state75_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state75_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state75_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state75_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state75_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state75_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state75_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state75_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state75_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state75_53_1 = reservoir_state[53] <<< 1;
wire signed [31:0] shifted_state75_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state75_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state75_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state75_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state75_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state75_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state75_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state75_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state75_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state75_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state75_88_5 = reservoir_state[88] <<< 5;
wire signed [31:0] shifted_state75_88_6 = reservoir_state[88] <<< 6;
wire signed [31:0] shifted_state75_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state75_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state75_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state75_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state75_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state75_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state75_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state75_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state75_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state75_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state75_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state75_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state75_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state75_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state75_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state75_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state75_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state75_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state75_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state75_108_4 = reservoir_state[108] <<< 4;
wire signed [31:0] shifted_state75_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state75_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state75_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state75_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state75_126_3 = reservoir_state[126] <<< 3;
wire signed [31:0] shifted_state75_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state75_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state75_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state75_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state75_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state75_134_2 = reservoir_state[134] <<< 2;
wire signed [31:0] shifted_state75_134_5 = reservoir_state[134] <<< 5;
wire signed [31:0] shifted_state75_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state75_146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state75_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state75_146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state75_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state75_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state75_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state75_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state75_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state75_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state75_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state75_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state75_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state75_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state75_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state75_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state75_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state75_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state75_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state75_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state75_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state75_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state75_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state75_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state76_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state76_1_1 = reservoir_state[1] <<< 1;
wire signed [31:0] shifted_state76_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state76_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state76_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state76_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state76_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state76_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state76_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state76_33_4 = reservoir_state[33] <<< 4;
wire signed [31:0] shifted_state76_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state76_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state76_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state76_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state76_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state76_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state76_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state76_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state76_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state76_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state76_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state76_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state76_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state76_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state76_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state76_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state76_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state76_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state76_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state76_74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state76_74_3 = reservoir_state[74] <<< 3;
wire signed [31:0] shifted_state76_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state76_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state76_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state76_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state76_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state76_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state76_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state76_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state76_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state76_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state76_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state76_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state76_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state76_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state76_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state76_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state76_154_0 = reservoir_state[154] <<< 0;
wire signed [31:0] shifted_state76_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state76_154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state76_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state76_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state76_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state76_159_0 = reservoir_state[159] <<< 0;
wire signed [31:0] shifted_state76_159_1 = reservoir_state[159] <<< 1;
wire signed [31:0] shifted_state76_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state76_159_5 = reservoir_state[159] <<< 5;
wire signed [31:0] shifted_state76_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state76_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state76_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state76_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state76_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state76_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state76_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state77_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state77_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state77_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state77_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state77_55_2 = reservoir_state[55] <<< 2;
wire signed [31:0] shifted_state77_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state77_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state77_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state77_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state77_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state77_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state77_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state77_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state77_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state77_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state77_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state77_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state77_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state77_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state77_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state77_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state77_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state77_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state77_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state77_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state77_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state77_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state77_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state77_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state77_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state77_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state77_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state77_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state77_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state77_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state77_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state77_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state77_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state77_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state77_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state78_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state78_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state78_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state78_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state78_30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state78_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state78_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state78_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state78_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state78_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state78_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state78_52_0 = reservoir_state[52] <<< 0;
wire signed [31:0] shifted_state78_52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state78_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state78_52_5 = reservoir_state[52] <<< 5;
wire signed [31:0] shifted_state78_52_6 = reservoir_state[52] <<< 6;
wire signed [31:0] shifted_state78_52_7 = reservoir_state[52] <<< 7;
wire signed [31:0] shifted_state78_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state78_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state78_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state78_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state78_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state78_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state78_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state78_90_1 = reservoir_state[90] <<< 1;
wire signed [31:0] shifted_state78_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state78_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state78_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state78_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state78_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state78_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state78_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state78_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state78_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state78_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state78_125_2 = reservoir_state[125] <<< 2;
wire signed [31:0] shifted_state78_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state78_128_2 = reservoir_state[128] <<< 2;
wire signed [31:0] shifted_state78_128_4 = reservoir_state[128] <<< 4;
wire signed [31:0] shifted_state78_128_5 = reservoir_state[128] <<< 5;
wire signed [31:0] shifted_state78_128_6 = reservoir_state[128] <<< 6;
wire signed [31:0] shifted_state78_128_7 = reservoir_state[128] <<< 7;
wire signed [31:0] shifted_state78_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state78_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state78_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state78_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state78_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state78_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state78_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state78_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state78_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state78_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state78_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state78_162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state78_162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state78_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state78_171_5 = reservoir_state[171] <<< 5;
wire signed [31:0] shifted_state78_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state78_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state78_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state78_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state78_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state78_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state79_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state79_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state79_12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state79_12_2 = reservoir_state[12] <<< 2;
wire signed [31:0] shifted_state79_12_4 = reservoir_state[12] <<< 4;
wire signed [31:0] shifted_state79_15_0 = reservoir_state[15] <<< 0;
wire signed [31:0] shifted_state79_15_3 = reservoir_state[15] <<< 3;
wire signed [31:0] shifted_state79_15_4 = reservoir_state[15] <<< 4;
wire signed [31:0] shifted_state79_15_5 = reservoir_state[15] <<< 5;
wire signed [31:0] shifted_state79_15_6 = reservoir_state[15] <<< 6;
wire signed [31:0] shifted_state79_15_7 = reservoir_state[15] <<< 7;
wire signed [31:0] shifted_state79_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state79_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state79_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state79_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state79_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state79_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state79_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state79_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state79_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state79_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state79_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state79_72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state79_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state79_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state79_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state79_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state79_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state79_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state79_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state79_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state79_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state79_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state79_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state79_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state79_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state79_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state79_108_4 = reservoir_state[108] <<< 4;
wire signed [31:0] shifted_state79_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state79_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state79_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state79_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state79_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state79_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state79_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state79_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state79_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state79_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state79_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state79_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state79_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state79_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state79_144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state79_144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state79_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state79_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state79_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state79_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state79_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state79_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state79_158_3 = reservoir_state[158] <<< 3;
wire signed [31:0] shifted_state79_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state79_158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state79_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state79_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state79_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state79_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state79_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state79_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state79_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state79_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state79_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state79_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state79_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state79_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state79_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state79_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state79_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state79_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state79_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state79_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state79_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state79_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state79_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state79_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state80_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state80_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state80_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state80_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state80_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state80_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state80_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state80_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state80_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state80_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state80_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state80_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state80_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state80_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state80_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state80_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state80_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state80_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state80_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state80_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state80_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state80_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state80_52_1 = reservoir_state[52] <<< 1;
wire signed [31:0] shifted_state80_52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state80_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state80_52_4 = reservoir_state[52] <<< 4;
wire signed [31:0] shifted_state80_52_6 = reservoir_state[52] <<< 6;
wire signed [31:0] shifted_state80_52_7 = reservoir_state[52] <<< 7;
wire signed [31:0] shifted_state80_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state80_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state80_57_3 = reservoir_state[57] <<< 3;
wire signed [31:0] shifted_state80_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state80_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state80_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state80_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state80_67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state80_67_3 = reservoir_state[67] <<< 3;
wire signed [31:0] shifted_state80_67_4 = reservoir_state[67] <<< 4;
wire signed [31:0] shifted_state80_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state80_67_6 = reservoir_state[67] <<< 6;
wire signed [31:0] shifted_state80_67_7 = reservoir_state[67] <<< 7;
wire signed [31:0] shifted_state80_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state80_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state80_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state80_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state80_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state80_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state80_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state80_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state80_92_1 = reservoir_state[92] <<< 1;
wire signed [31:0] shifted_state80_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state80_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state80_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state80_94_2 = reservoir_state[94] <<< 2;
wire signed [31:0] shifted_state80_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state80_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state80_115_3 = reservoir_state[115] <<< 3;
wire signed [31:0] shifted_state80_115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state80_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state80_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state80_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state80_153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state80_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state80_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state80_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state80_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state80_158_0 = reservoir_state[158] <<< 0;
wire signed [31:0] shifted_state80_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state80_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state80_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state80_158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state80_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state80_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state80_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state80_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state80_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state80_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state80_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state80_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state80_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state80_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state80_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state80_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state80_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state80_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state80_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state80_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state80_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state80_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state80_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state80_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state80_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state80_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state80_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state80_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state80_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state81_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state81_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state81_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state81_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state81_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state81_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state81_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state81_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state81_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state81_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state81_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state81_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state81_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state81_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state81_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state81_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state81_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state81_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state81_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state81_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state81_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state81_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state81_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state81_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state81_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state81_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state81_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state81_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state81_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state81_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state81_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state81_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state81_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state81_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state81_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state81_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state81_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state81_56_5 = reservoir_state[56] <<< 5;
wire signed [31:0] shifted_state81_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state81_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state81_58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state81_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state81_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state81_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state81_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state81_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state81_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state81_64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state81_64_6 = reservoir_state[64] <<< 6;
wire signed [31:0] shifted_state81_64_7 = reservoir_state[64] <<< 7;
wire signed [31:0] shifted_state81_74_3 = reservoir_state[74] <<< 3;
wire signed [31:0] shifted_state81_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state81_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state81_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state81_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state81_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state81_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state81_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state81_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state81_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state81_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state81_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state81_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state81_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state81_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state81_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state81_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state81_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state81_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state81_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state81_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state81_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state81_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state81_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state81_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state81_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state81_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state81_146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state81_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state81_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state81_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state81_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state81_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state81_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state81_171_6 = reservoir_state[171] <<< 6;
wire signed [31:0] shifted_state81_171_7 = reservoir_state[171] <<< 7;
wire signed [31:0] shifted_state81_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state81_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state82_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state82_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state82_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state82_8_1 = reservoir_state[8] <<< 1;
wire signed [31:0] shifted_state82_12_0 = reservoir_state[12] <<< 0;
wire signed [31:0] shifted_state82_12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state82_12_3 = reservoir_state[12] <<< 3;
wire signed [31:0] shifted_state82_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state82_15_3 = reservoir_state[15] <<< 3;
wire signed [31:0] shifted_state82_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state82_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state82_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state82_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state82_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state82_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state82_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state82_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state82_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state82_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state82_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state82_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state82_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state82_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state82_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state82_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state82_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state82_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state82_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state82_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state82_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state82_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state82_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state82_91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state82_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state82_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state82_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state82_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state82_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state82_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state82_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state82_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state82_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state82_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state82_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state82_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state82_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state82_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state82_136_2 = reservoir_state[136] <<< 2;
wire signed [31:0] shifted_state82_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state82_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state82_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state82_146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state82_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state82_146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state82_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state82_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state82_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state82_149_1 = reservoir_state[149] <<< 1;
wire signed [31:0] shifted_state82_149_2 = reservoir_state[149] <<< 2;
wire signed [31:0] shifted_state82_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state82_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state82_149_5 = reservoir_state[149] <<< 5;
wire signed [31:0] shifted_state82_149_7 = reservoir_state[149] <<< 7;
wire signed [31:0] shifted_state82_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state82_154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state82_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state82_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state82_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state82_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state82_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state82_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state82_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state82_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state82_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state82_167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state82_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state82_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state82_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state82_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state82_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state82_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state82_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state82_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state82_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state82_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state82_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state82_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state82_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state83_8_1 = reservoir_state[8] <<< 1;
wire signed [31:0] shifted_state83_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state83_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state83_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state83_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state83_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state83_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state83_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state83_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state83_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state83_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state83_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state83_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state83_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state83_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state83_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state83_36_4 = reservoir_state[36] <<< 4;
wire signed [31:0] shifted_state83_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state83_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state83_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state83_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state83_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state83_47_4 = reservoir_state[47] <<< 4;
wire signed [31:0] shifted_state83_47_5 = reservoir_state[47] <<< 5;
wire signed [31:0] shifted_state83_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state83_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state83_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state83_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state83_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state83_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state83_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state83_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state83_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state83_75_2 = reservoir_state[75] <<< 2;
wire signed [31:0] shifted_state83_75_3 = reservoir_state[75] <<< 3;
wire signed [31:0] shifted_state83_75_4 = reservoir_state[75] <<< 4;
wire signed [31:0] shifted_state83_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state83_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state83_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state83_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state83_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state83_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state83_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state83_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state83_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state83_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state83_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state83_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state83_108_4 = reservoir_state[108] <<< 4;
wire signed [31:0] shifted_state83_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state83_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state83_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state83_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state83_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state83_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state83_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state83_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state83_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state83_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state83_156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state84_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state84_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state84_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state84_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state84_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state84_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state84_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state84_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state84_70_4 = reservoir_state[70] <<< 4;
wire signed [31:0] shifted_state84_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state84_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state84_74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state84_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state84_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state84_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state84_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state84_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state84_79_5 = reservoir_state[79] <<< 5;
wire signed [31:0] shifted_state84_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state84_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state84_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state84_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state84_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state84_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state84_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state84_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state84_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state84_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state84_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state84_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state84_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state84_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state84_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state84_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state84_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state84_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state84_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state84_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state84_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state84_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state84_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state84_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state84_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state84_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state84_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state84_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state84_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state84_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state84_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state84_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state84_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state84_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state84_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state84_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state84_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state84_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state84_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state84_194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state84_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state84_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state84_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state85_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state85_2_3 = reservoir_state[2] <<< 3;
wire signed [31:0] shifted_state85_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state85_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state85_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state85_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state85_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state85_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state85_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state85_13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state85_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state85_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state85_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state85_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state85_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state85_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state85_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state85_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state85_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state85_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state85_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state85_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state85_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state85_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state85_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state85_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state85_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state85_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state85_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state85_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state85_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state85_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state85_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state85_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state85_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state85_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state85_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state85_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state85_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state85_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state85_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state85_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state85_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state85_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state85_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state85_75_5 = reservoir_state[75] <<< 5;
wire signed [31:0] shifted_state85_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state85_81_2 = reservoir_state[81] <<< 2;
wire signed [31:0] shifted_state85_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state85_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state85_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state85_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state85_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state85_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state85_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state85_88_5 = reservoir_state[88] <<< 5;
wire signed [31:0] shifted_state85_88_6 = reservoir_state[88] <<< 6;
wire signed [31:0] shifted_state85_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state85_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state85_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state85_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state85_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state85_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state85_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state85_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state85_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state85_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state85_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state85_161_0 = reservoir_state[161] <<< 0;
wire signed [31:0] shifted_state85_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state85_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state85_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state85_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state85_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state85_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state85_176_0 = reservoir_state[176] <<< 0;
wire signed [31:0] shifted_state85_176_4 = reservoir_state[176] <<< 4;
wire signed [31:0] shifted_state85_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state85_181_1 = reservoir_state[181] <<< 1;
wire signed [31:0] shifted_state85_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state85_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state85_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state85_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state85_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state85_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state85_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state85_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state85_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state85_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state85_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state85_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state85_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state85_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state85_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state85_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state85_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state85_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state85_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state85_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state85_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state85_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state85_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state85_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state85_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state85_196_6 = reservoir_state[196] <<< 6;
wire signed [31:0] shifted_state86_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state86_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state86_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state86_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state86_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state86_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state86_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state86_9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state86_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state86_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state86_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state86_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state86_18_3 = reservoir_state[18] <<< 3;
wire signed [31:0] shifted_state86_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state86_40_5 = reservoir_state[40] <<< 5;
wire signed [31:0] shifted_state86_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state86_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state86_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state86_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state86_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state86_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state86_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state86_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state86_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state86_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state86_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state86_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state86_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state86_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state86_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state86_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state86_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state86_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state86_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state86_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state86_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state86_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state86_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state86_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state86_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state86_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state86_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state86_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state86_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state86_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state86_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state86_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state86_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state86_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state86_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state86_88_6 = reservoir_state[88] <<< 6;
wire signed [31:0] shifted_state86_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state86_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state86_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state86_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state86_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state86_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state86_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state86_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state86_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state86_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state86_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state86_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state86_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state86_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state86_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state86_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state86_118_3 = reservoir_state[118] <<< 3;
wire signed [31:0] shifted_state86_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state86_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state86_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state86_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state86_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state86_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state86_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state86_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state86_137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state86_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state86_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state86_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state86_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state86_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state86_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state86_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state86_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state86_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state86_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state86_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state86_153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state86_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state86_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state86_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state86_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state86_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state86_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state86_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state86_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state86_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state86_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state86_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state86_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state86_169_2 = reservoir_state[169] <<< 2;
wire signed [31:0] shifted_state86_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state86_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state86_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state86_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state86_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state86_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state86_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state86_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state86_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state86_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state86_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state86_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state86_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state86_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state86_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state86_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state86_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state86_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state86_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state86_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state86_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state86_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state86_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state86_199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state86_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state86_199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state87_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state87_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state87_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state87_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state87_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state87_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state87_12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state87_12_2 = reservoir_state[12] <<< 2;
wire signed [31:0] shifted_state87_12_6 = reservoir_state[12] <<< 6;
wire signed [31:0] shifted_state87_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state87_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state87_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state87_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state87_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state87_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state87_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state87_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state87_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state87_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state87_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state87_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state87_40_2 = reservoir_state[40] <<< 2;
wire signed [31:0] shifted_state87_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state87_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state87_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state87_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state87_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state87_48_5 = reservoir_state[48] <<< 5;
wire signed [31:0] shifted_state87_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state87_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state87_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state87_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state87_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state87_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state87_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state87_60_4 = reservoir_state[60] <<< 4;
wire signed [31:0] shifted_state87_67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state87_67_1 = reservoir_state[67] <<< 1;
wire signed [31:0] shifted_state87_67_2 = reservoir_state[67] <<< 2;
wire signed [31:0] shifted_state87_67_3 = reservoir_state[67] <<< 3;
wire signed [31:0] shifted_state87_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state87_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state87_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state87_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state87_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state87_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state87_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state87_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state87_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state87_101_2 = reservoir_state[101] <<< 2;
wire signed [31:0] shifted_state87_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state87_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state87_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state87_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state87_103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state87_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state87_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state87_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state87_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state87_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state87_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state87_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state87_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state87_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state87_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state87_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state87_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state87_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state87_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state87_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state87_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state87_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state87_131_4 = reservoir_state[131] <<< 4;
wire signed [31:0] shifted_state87_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state87_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state87_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state87_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state87_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state87_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state87_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state87_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state87_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state87_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state87_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state87_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state87_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state87_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state87_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state87_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state87_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state87_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state87_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state87_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state87_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state88_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state88_1_1 = reservoir_state[1] <<< 1;
wire signed [31:0] shifted_state88_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state88_1_3 = reservoir_state[1] <<< 3;
wire signed [31:0] shifted_state88_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state88_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state88_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state88_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state88_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state88_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state88_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state88_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state88_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state88_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state88_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state88_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state88_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state88_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state88_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state88_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state88_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state88_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state88_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state88_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state88_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state88_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state88_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state88_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state88_74_3 = reservoir_state[74] <<< 3;
wire signed [31:0] shifted_state88_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state88_92_1 = reservoir_state[92] <<< 1;
wire signed [31:0] shifted_state88_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state88_92_4 = reservoir_state[92] <<< 4;
wire signed [31:0] shifted_state88_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state88_103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state88_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state88_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state88_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state88_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state88_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state88_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state88_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state88_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state88_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state88_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state88_154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state88_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state88_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state88_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state88_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state88_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state88_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state88_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state88_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state88_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state88_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state88_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state88_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state88_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state88_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state88_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state88_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state88_197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state88_197_4 = reservoir_state[197] <<< 4;
wire signed [31:0] shifted_state88_197_5 = reservoir_state[197] <<< 5;
wire signed [31:0] shifted_state88_197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state88_197_7 = reservoir_state[197] <<< 7;
wire signed [31:0] shifted_state89_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state89_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state89_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state89_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state89_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state89_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state89_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state89_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state89_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state89_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state89_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state89_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state89_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state89_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state89_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state89_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state89_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state89_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state89_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state89_50_4 = reservoir_state[50] <<< 4;
wire signed [31:0] shifted_state89_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state89_58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state89_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state89_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state89_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state89_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state89_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state89_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state89_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state89_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state89_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state89_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state89_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state89_74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state89_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state89_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state89_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state89_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state89_79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state89_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state89_79_5 = reservoir_state[79] <<< 5;
wire signed [31:0] shifted_state89_79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state89_79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state89_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state89_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state89_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state89_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state89_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state89_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state89_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state89_122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state89_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state89_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state89_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state89_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state89_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state89_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state89_134_0 = reservoir_state[134] <<< 0;
wire signed [31:0] shifted_state89_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state89_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state89_134_4 = reservoir_state[134] <<< 4;
wire signed [31:0] shifted_state89_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state89_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state89_144_0 = reservoir_state[144] <<< 0;
wire signed [31:0] shifted_state89_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state89_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state89_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state89_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state89_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state89_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state89_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state89_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state89_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state89_156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state89_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state89_176_2 = reservoir_state[176] <<< 2;
wire signed [31:0] shifted_state89_176_3 = reservoir_state[176] <<< 3;
wire signed [31:0] shifted_state89_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state89_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state89_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state89_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state89_181_1 = reservoir_state[181] <<< 1;
wire signed [31:0] shifted_state89_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state89_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state89_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state89_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state89_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state89_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state89_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state89_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state89_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state89_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state89_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state89_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state89_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state89_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state89_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state89_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state89_189_6 = reservoir_state[189] <<< 6;
wire signed [31:0] shifted_state89_189_7 = reservoir_state[189] <<< 7;
wire signed [31:0] shifted_state90_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state90_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state90_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state90_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state90_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state90_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state90_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state90_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state90_6_3 = reservoir_state[6] <<< 3;
wire signed [31:0] shifted_state90_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state90_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state90_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state90_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state90_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state90_19_1 = reservoir_state[19] <<< 1;
wire signed [31:0] shifted_state90_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state90_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state90_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state90_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state90_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state90_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state90_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state90_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state90_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state90_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state90_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state90_69_1 = reservoir_state[69] <<< 1;
wire signed [31:0] shifted_state90_69_2 = reservoir_state[69] <<< 2;
wire signed [31:0] shifted_state90_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state90_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state90_69_6 = reservoir_state[69] <<< 6;
wire signed [31:0] shifted_state90_69_7 = reservoir_state[69] <<< 7;
wire signed [31:0] shifted_state90_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state90_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state90_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state90_114_1 = reservoir_state[114] <<< 1;
wire signed [31:0] shifted_state90_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state90_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state90_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state90_117_5 = reservoir_state[117] <<< 5;
wire signed [31:0] shifted_state90_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state90_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state90_122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state90_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state90_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state90_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state90_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state90_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state90_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state90_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state90_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state90_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state90_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state90_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state90_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state90_167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state90_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state90_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state90_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state90_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state91_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state91_3_1 = reservoir_state[3] <<< 1;
wire signed [31:0] shifted_state91_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state91_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state91_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state91_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state91_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state91_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state91_29_2 = reservoir_state[29] <<< 2;
wire signed [31:0] shifted_state91_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state91_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state91_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state91_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state91_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state91_56_0 = reservoir_state[56] <<< 0;
wire signed [31:0] shifted_state91_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state91_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state91_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state91_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state91_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state91_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state91_64_4 = reservoir_state[64] <<< 4;
wire signed [31:0] shifted_state91_64_6 = reservoir_state[64] <<< 6;
wire signed [31:0] shifted_state91_64_7 = reservoir_state[64] <<< 7;
wire signed [31:0] shifted_state91_73_3 = reservoir_state[73] <<< 3;
wire signed [31:0] shifted_state91_73_5 = reservoir_state[73] <<< 5;
wire signed [31:0] shifted_state91_73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state91_73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state91_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state91_87_1 = reservoir_state[87] <<< 1;
wire signed [31:0] shifted_state91_87_3 = reservoir_state[87] <<< 3;
wire signed [31:0] shifted_state91_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state91_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state91_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state91_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state91_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state91_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state91_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state91_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state91_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state91_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state91_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state91_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state91_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state91_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state91_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state91_103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state91_103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state91_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state91_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state91_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state91_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state91_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state91_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state91_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state91_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state91_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state91_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state91_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state91_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state91_142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state91_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state91_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state91_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state91_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state91_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state91_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state91_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state91_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state91_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state91_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state91_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state91_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state91_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state91_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state91_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state91_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state91_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state91_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state91_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state91_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state91_194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state91_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state91_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state91_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state91_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state91_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state92_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state92_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state92_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state92_18_3 = reservoir_state[18] <<< 3;
wire signed [31:0] shifted_state92_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state92_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state92_39_0 = reservoir_state[39] <<< 0;
wire signed [31:0] shifted_state92_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state92_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state92_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state92_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state92_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state92_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state92_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state92_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state92_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state92_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state92_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state92_84_2 = reservoir_state[84] <<< 2;
wire signed [31:0] shifted_state92_84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state92_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state92_84_5 = reservoir_state[84] <<< 5;
wire signed [31:0] shifted_state92_84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state92_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state92_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state92_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state92_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state92_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state92_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state92_103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state92_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state92_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state92_119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state92_119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state92_119_3 = reservoir_state[119] <<< 3;
wire signed [31:0] shifted_state92_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state92_119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state92_119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state92_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state92_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state92_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state92_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state92_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state92_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state92_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state92_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state92_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state92_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state92_137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state92_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state92_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state92_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state92_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state92_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state92_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state92_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state92_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state92_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state92_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state92_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state92_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state92_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state92_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state92_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state92_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state92_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state92_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state92_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state92_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state93_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state93_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state93_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state93_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state93_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state93_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state93_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state93_27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state93_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state93_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state93_27_6 = reservoir_state[27] <<< 6;
wire signed [31:0] shifted_state93_27_7 = reservoir_state[27] <<< 7;
wire signed [31:0] shifted_state93_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state93_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state93_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state93_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state93_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state93_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state93_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state93_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state93_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state93_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state93_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state93_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state93_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state93_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state93_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state93_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state93_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state93_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state93_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state93_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state93_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state93_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state93_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state93_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state93_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state93_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state93_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state93_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state93_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state93_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state93_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state93_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state93_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state93_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state93_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state93_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state93_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state93_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state93_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state93_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state93_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state93_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state93_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state93_112_3 = reservoir_state[112] <<< 3;
wire signed [31:0] shifted_state93_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state93_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state93_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state93_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state93_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state93_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state93_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state93_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state93_143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state93_143_2 = reservoir_state[143] <<< 2;
wire signed [31:0] shifted_state93_143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state93_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state93_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state93_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state93_149_2 = reservoir_state[149] <<< 2;
wire signed [31:0] shifted_state93_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state93_149_5 = reservoir_state[149] <<< 5;
wire signed [31:0] shifted_state93_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state93_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state93_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state93_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state93_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state93_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state93_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state93_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state93_151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state93_151_4 = reservoir_state[151] <<< 4;
wire signed [31:0] shifted_state93_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state93_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state93_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state93_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state93_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state93_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state93_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state93_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state93_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state93_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state93_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state93_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state93_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state93_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state93_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state93_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state93_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state93_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state93_185_2 = reservoir_state[185] <<< 2;
wire signed [31:0] shifted_state94_2_0 = reservoir_state[2] <<< 0;
wire signed [31:0] shifted_state94_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state94_2_3 = reservoir_state[2] <<< 3;
wire signed [31:0] shifted_state94_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state94_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state94_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state94_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state94_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state94_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state94_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state94_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state94_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state94_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state94_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state94_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state94_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state94_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state94_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state94_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state94_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state94_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state94_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state94_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state94_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state94_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state94_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state94_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state94_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state94_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state94_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state94_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state94_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state94_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state94_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state94_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state94_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state94_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state94_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state94_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state94_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state94_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state94_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state94_84_5 = reservoir_state[84] <<< 5;
wire signed [31:0] shifted_state94_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state94_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state94_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state94_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state94_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state94_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state94_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state94_102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state94_102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state94_102_7 = reservoir_state[102] <<< 7;
wire signed [31:0] shifted_state94_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state94_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state94_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state94_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state94_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state94_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state94_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state94_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state94_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state94_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state94_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state94_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state94_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state94_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state94_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state94_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state94_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state94_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state94_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state94_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state94_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state94_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state94_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state94_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state94_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state94_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state95_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state95_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state95_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state95_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state95_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state95_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state95_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state95_30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state95_30_5 = reservoir_state[30] <<< 5;
wire signed [31:0] shifted_state95_30_6 = reservoir_state[30] <<< 6;
wire signed [31:0] shifted_state95_30_7 = reservoir_state[30] <<< 7;
wire signed [31:0] shifted_state95_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state95_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state95_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state95_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state95_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state95_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state95_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state95_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state95_73_2 = reservoir_state[73] <<< 2;
wire signed [31:0] shifted_state95_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state95_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state95_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state95_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state95_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state95_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state95_98_5 = reservoir_state[98] <<< 5;
wire signed [31:0] shifted_state95_98_6 = reservoir_state[98] <<< 6;
wire signed [31:0] shifted_state95_98_7 = reservoir_state[98] <<< 7;
wire signed [31:0] shifted_state95_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state95_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state95_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state95_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state95_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state95_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state95_117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state95_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state95_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state95_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state95_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state95_147_1 = reservoir_state[147] <<< 1;
wire signed [31:0] shifted_state95_147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state95_147_3 = reservoir_state[147] <<< 3;
wire signed [31:0] shifted_state95_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state95_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state95_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state95_149_5 = reservoir_state[149] <<< 5;
wire signed [31:0] shifted_state95_159_0 = reservoir_state[159] <<< 0;
wire signed [31:0] shifted_state95_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state95_159_4 = reservoir_state[159] <<< 4;
wire signed [31:0] shifted_state95_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state95_161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state95_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state95_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state95_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state95_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state95_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state95_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state95_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state95_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state95_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state95_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state95_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state95_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state95_171_0 = reservoir_state[171] <<< 0;
wire signed [31:0] shifted_state95_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state95_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state95_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state95_176_3 = reservoir_state[176] <<< 3;
wire signed [31:0] shifted_state95_176_5 = reservoir_state[176] <<< 5;
wire signed [31:0] shifted_state95_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state95_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state95_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state95_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state95_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state95_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state95_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state95_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state96_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state96_3_1 = reservoir_state[3] <<< 1;
wire signed [31:0] shifted_state96_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state96_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state96_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state96_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state96_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state96_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state96_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state96_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state96_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state96_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state96_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state96_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state96_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state96_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state96_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state96_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state96_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state96_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state96_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state96_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state96_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state96_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state96_48_5 = reservoir_state[48] <<< 5;
wire signed [31:0] shifted_state96_48_6 = reservoir_state[48] <<< 6;
wire signed [31:0] shifted_state96_48_7 = reservoir_state[48] <<< 7;
wire signed [31:0] shifted_state96_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state96_49_1 = reservoir_state[49] <<< 1;
wire signed [31:0] shifted_state96_49_4 = reservoir_state[49] <<< 4;
wire signed [31:0] shifted_state96_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state96_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state96_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state96_52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state96_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state96_52_5 = reservoir_state[52] <<< 5;
wire signed [31:0] shifted_state96_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state96_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state96_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state96_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state96_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state96_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state96_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state96_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state96_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state96_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state96_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state96_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state96_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state96_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state96_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state96_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state96_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state96_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state96_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state96_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state96_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state96_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state96_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state96_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state96_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state96_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state96_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state96_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state96_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state96_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state96_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state96_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state96_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state96_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state96_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state96_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state96_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state96_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state96_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state96_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state96_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state96_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state97_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state97_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state97_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state97_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state97_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state97_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state97_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state97_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state97_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state97_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state97_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state97_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state97_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state97_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state97_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state97_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state97_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state97_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state97_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state97_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state97_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state97_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state97_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state97_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state97_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state97_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state97_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state97_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state97_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state97_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state97_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state97_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state97_135_3 = reservoir_state[135] <<< 3;
wire signed [31:0] shifted_state97_135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state97_135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state97_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state97_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state97_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state97_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state97_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state97_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state97_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state97_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state97_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state97_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state97_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state97_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state97_167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state97_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state97_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state97_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state97_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state97_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state97_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state97_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state97_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state97_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state98_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state98_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state98_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state98_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state98_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state98_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state98_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state98_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state98_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state98_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state98_43_1 = reservoir_state[43] <<< 1;
wire signed [31:0] shifted_state98_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state98_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state98_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state98_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state98_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state98_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state98_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state98_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state98_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state98_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state98_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state98_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state98_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state98_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state98_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state98_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state98_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state98_75_1 = reservoir_state[75] <<< 1;
wire signed [31:0] shifted_state98_75_2 = reservoir_state[75] <<< 2;
wire signed [31:0] shifted_state98_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state98_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state98_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state98_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state98_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state98_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state98_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state98_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state98_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state98_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state98_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state98_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state98_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state98_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state98_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state98_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state98_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state98_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state98_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state98_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state98_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state98_102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state98_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state98_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state98_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state98_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state98_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state98_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state98_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state98_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state98_115_3 = reservoir_state[115] <<< 3;
wire signed [31:0] shifted_state98_115_4 = reservoir_state[115] <<< 4;
wire signed [31:0] shifted_state98_115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state98_115_6 = reservoir_state[115] <<< 6;
wire signed [31:0] shifted_state98_115_7 = reservoir_state[115] <<< 7;
wire signed [31:0] shifted_state98_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state98_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state98_119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state98_119_2 = reservoir_state[119] <<< 2;
wire signed [31:0] shifted_state98_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state98_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state98_119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state98_119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state98_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state98_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state98_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state98_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state98_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state98_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state98_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state98_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state98_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state98_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state98_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state98_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state98_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state98_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state98_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state98_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state98_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state98_196_0 = reservoir_state[196] <<< 0;
wire signed [31:0] shifted_state98_196_1 = reservoir_state[196] <<< 1;
wire signed [31:0] shifted_state98_196_3 = reservoir_state[196] <<< 3;
wire signed [31:0] shifted_state98_196_4 = reservoir_state[196] <<< 4;
wire signed [31:0] shifted_state98_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state98_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state98_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state98_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state98_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state99_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state99_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state99_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state99_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state99_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state99_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state99_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state99_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state99_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state99_2_3 = reservoir_state[2] <<< 3;
wire signed [31:0] shifted_state99_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state99_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state99_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state99_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state99_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state99_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state99_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state99_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state99_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state99_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state99_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state99_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state99_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state99_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state99_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state99_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state99_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state99_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state99_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state99_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state99_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state99_56_5 = reservoir_state[56] <<< 5;
wire signed [31:0] shifted_state99_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state99_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state99_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state99_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state99_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state99_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state99_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state99_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state99_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state99_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state99_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state99_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state99_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state99_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state99_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state99_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state99_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state99_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state99_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state99_90_4 = reservoir_state[90] <<< 4;
wire signed [31:0] shifted_state99_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state99_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state99_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state99_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state99_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state99_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state99_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state99_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state99_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state99_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state99_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state99_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state99_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state99_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state99_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state99_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state99_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state99_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state99_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state99_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state99_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state99_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state99_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state99_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state99_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state99_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state99_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state99_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state99_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state99_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state99_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state99_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state99_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state99_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state99_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state99_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state99_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state99_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state99_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state99_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state99_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state99_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state99_142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state99_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state99_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state99_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state99_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state99_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state99_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state99_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state99_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state99_156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state99_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state99_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state99_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state99_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state99_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state99_197_2 = reservoir_state[197] <<< 2;
wire signed [31:0] shifted_state99_197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state99_197_4 = reservoir_state[197] <<< 4;
wire signed [31:0] shifted_state99_197_5 = reservoir_state[197] <<< 5;
wire signed [31:0] shifted_state100_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state100_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state100_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state100_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state100_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state100_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state100_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state100_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state100_29_5 = reservoir_state[29] <<< 5;
wire signed [31:0] shifted_state100_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state100_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state100_39_0 = reservoir_state[39] <<< 0;
wire signed [31:0] shifted_state100_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state100_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state100_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state100_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state100_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state100_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state100_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state100_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state100_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state100_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state100_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state100_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state100_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state100_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state100_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state100_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state100_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state100_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state100_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state100_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state100_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state100_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state100_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state100_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state100_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state100_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state100_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state100_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state100_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state100_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state100_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state100_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state100_120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state100_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state100_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state100_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state100_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state100_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state100_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state100_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state100_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state100_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state100_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state100_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state100_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state100_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state100_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state100_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state100_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state100_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state100_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state100_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state100_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state100_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state100_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state100_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state100_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state100_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state100_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state100_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state100_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state100_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state100_199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state100_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state100_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state101_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state101_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state101_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state101_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state101_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state101_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state101_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state101_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state101_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state101_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state101_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state101_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state101_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state101_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state101_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state101_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state101_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state101_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state101_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state101_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state101_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state101_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state101_56_5 = reservoir_state[56] <<< 5;
wire signed [31:0] shifted_state101_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state101_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state101_81_2 = reservoir_state[81] <<< 2;
wire signed [31:0] shifted_state101_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state101_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state101_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state101_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state101_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state101_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state101_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state101_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state101_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state101_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state101_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state101_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state101_92_1 = reservoir_state[92] <<< 1;
wire signed [31:0] shifted_state101_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state101_92_6 = reservoir_state[92] <<< 6;
wire signed [31:0] shifted_state101_92_7 = reservoir_state[92] <<< 7;
wire signed [31:0] shifted_state101_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state101_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state101_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state101_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state101_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state101_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state101_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state101_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state101_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state101_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state101_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state101_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state101_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state101_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state101_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state101_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state101_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state101_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state101_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state101_149_6 = reservoir_state[149] <<< 6;
wire signed [31:0] shifted_state101_149_7 = reservoir_state[149] <<< 7;
wire signed [31:0] shifted_state101_157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state101_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state101_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state101_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state101_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state101_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state101_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state101_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state101_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state101_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state102_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state102_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state102_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state102_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state102_16_3 = reservoir_state[16] <<< 3;
wire signed [31:0] shifted_state102_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state102_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state102_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state102_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state102_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state102_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state102_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state102_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state102_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state102_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state102_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state102_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state102_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state102_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state102_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state102_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state102_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state102_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state102_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state102_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state102_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state102_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state102_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state102_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state102_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state102_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state102_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state102_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state102_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state102_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state102_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state102_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state102_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state102_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state102_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state102_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state102_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state102_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state102_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state102_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state102_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state102_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state102_102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state102_102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state102_102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state102_102_7 = reservoir_state[102] <<< 7;
wire signed [31:0] shifted_state102_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state102_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state102_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state102_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state102_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state102_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state102_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state102_120_2 = reservoir_state[120] <<< 2;
wire signed [31:0] shifted_state102_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state102_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state102_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state102_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state102_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state102_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state102_135_2 = reservoir_state[135] <<< 2;
wire signed [31:0] shifted_state102_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state102_135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state102_135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state102_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state102_146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state102_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state102_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state102_146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state102_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state102_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state102_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state102_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state102_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state102_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state102_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state102_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state102_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state102_171_6 = reservoir_state[171] <<< 6;
wire signed [31:0] shifted_state102_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state102_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state102_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state103_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state103_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state103_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state103_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state103_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state103_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state103_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state103_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state103_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state103_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state103_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state103_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state103_16_3 = reservoir_state[16] <<< 3;
wire signed [31:0] shifted_state103_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state103_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state103_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state103_29_5 = reservoir_state[29] <<< 5;
wire signed [31:0] shifted_state103_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state103_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state103_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state103_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state103_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state103_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state103_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state103_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state103_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state103_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state103_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state103_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state103_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state103_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state103_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state103_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state103_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state103_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state103_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state103_47_4 = reservoir_state[47] <<< 4;
wire signed [31:0] shifted_state103_47_5 = reservoir_state[47] <<< 5;
wire signed [31:0] shifted_state103_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state103_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state103_50_4 = reservoir_state[50] <<< 4;
wire signed [31:0] shifted_state103_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state103_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state103_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state103_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state103_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state103_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state103_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state103_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state103_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state103_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state103_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state103_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state103_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state103_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state103_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state103_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state103_73_2 = reservoir_state[73] <<< 2;
wire signed [31:0] shifted_state103_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state103_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state103_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state103_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state103_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state103_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state103_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state103_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state103_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state103_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state103_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state103_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state103_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state103_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state103_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state103_112_3 = reservoir_state[112] <<< 3;
wire signed [31:0] shifted_state103_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state103_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state103_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state103_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state103_136_2 = reservoir_state[136] <<< 2;
wire signed [31:0] shifted_state103_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state103_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state103_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state103_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state103_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state103_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state104_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state104_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state104_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state104_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state104_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state104_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state104_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state104_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state104_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state104_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state104_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state104_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state104_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state104_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state104_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state104_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state104_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state104_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state104_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state104_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state104_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state104_90_0 = reservoir_state[90] <<< 0;
wire signed [31:0] shifted_state104_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state104_90_4 = reservoir_state[90] <<< 4;
wire signed [31:0] shifted_state104_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state104_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state104_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state104_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state104_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state104_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state104_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state104_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state104_136_2 = reservoir_state[136] <<< 2;
wire signed [31:0] shifted_state104_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state104_140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state104_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state104_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state104_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state104_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state104_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state104_159_2 = reservoir_state[159] <<< 2;
wire signed [31:0] shifted_state104_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state104_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state104_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state104_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state104_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state104_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state104_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state104_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state104_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state104_171_5 = reservoir_state[171] <<< 5;
wire signed [31:0] shifted_state104_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state104_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state104_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state104_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state104_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state104_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state104_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state105_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state105_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state105_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state105_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state105_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state105_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state105_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state105_2_3 = reservoir_state[2] <<< 3;
wire signed [31:0] shifted_state105_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state105_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state105_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state105_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state105_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state105_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state105_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state105_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state105_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state105_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state105_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state105_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state105_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state105_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state105_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state105_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state105_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state105_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state105_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state105_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state105_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state105_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state105_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state105_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state105_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state105_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state105_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state105_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state105_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state105_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state105_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state105_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state105_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state105_70_0 = reservoir_state[70] <<< 0;
wire signed [31:0] shifted_state105_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state105_70_2 = reservoir_state[70] <<< 2;
wire signed [31:0] shifted_state105_70_4 = reservoir_state[70] <<< 4;
wire signed [31:0] shifted_state105_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state105_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state105_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state105_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state105_87_2 = reservoir_state[87] <<< 2;
wire signed [31:0] shifted_state105_87_3 = reservoir_state[87] <<< 3;
wire signed [31:0] shifted_state105_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state105_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state105_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state105_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state105_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state105_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state105_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state105_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state105_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state105_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state105_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state105_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state105_102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state105_102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state105_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state105_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state105_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state105_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state105_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state105_110_3 = reservoir_state[110] <<< 3;
wire signed [31:0] shifted_state105_110_4 = reservoir_state[110] <<< 4;
wire signed [31:0] shifted_state105_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state105_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state105_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state105_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state105_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state105_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state105_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state105_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state105_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state105_118_3 = reservoir_state[118] <<< 3;
wire signed [31:0] shifted_state105_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state105_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state105_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state105_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state105_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state105_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state105_120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state105_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state105_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state105_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state105_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state105_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state105_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state105_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state105_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state105_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state105_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state105_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state105_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state105_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state105_154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state105_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state105_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state105_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state105_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state105_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state105_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state105_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state105_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state106_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state106_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state106_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state106_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state106_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state106_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state106_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state106_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state106_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state106_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state106_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state106_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state106_23_4 = reservoir_state[23] <<< 4;
wire signed [31:0] shifted_state106_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state106_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state106_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state106_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state106_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state106_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state106_52_1 = reservoir_state[52] <<< 1;
wire signed [31:0] shifted_state106_52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state106_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state106_52_5 = reservoir_state[52] <<< 5;
wire signed [31:0] shifted_state106_52_6 = reservoir_state[52] <<< 6;
wire signed [31:0] shifted_state106_52_7 = reservoir_state[52] <<< 7;
wire signed [31:0] shifted_state106_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state106_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state106_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state106_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state106_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state106_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state106_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state106_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state106_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state106_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state106_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state106_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state106_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state106_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state106_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state106_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state106_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state106_114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state106_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state106_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state106_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state106_120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state106_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state106_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state106_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state106_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state106_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state106_144_0 = reservoir_state[144] <<< 0;
wire signed [31:0] shifted_state106_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state106_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state106_144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state106_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state106_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state106_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state106_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state106_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state106_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state106_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state106_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state106_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state106_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state106_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state106_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state106_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state106_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state106_199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state107_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state107_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state107_5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state107_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state107_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state107_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state107_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state107_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state107_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state107_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state107_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state107_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state107_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state107_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state107_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state107_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state107_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state107_48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state107_48_5 = reservoir_state[48] <<< 5;
wire signed [31:0] shifted_state107_48_7 = reservoir_state[48] <<< 7;
wire signed [31:0] shifted_state107_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state107_49_3 = reservoir_state[49] <<< 3;
wire signed [31:0] shifted_state107_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state107_75_3 = reservoir_state[75] <<< 3;
wire signed [31:0] shifted_state107_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state107_82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state107_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state107_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state107_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state107_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state107_120_2 = reservoir_state[120] <<< 2;
wire signed [31:0] shifted_state107_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state107_120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state107_120_5 = reservoir_state[120] <<< 5;
wire signed [31:0] shifted_state107_120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state107_120_7 = reservoir_state[120] <<< 7;
wire signed [31:0] shifted_state107_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state107_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state107_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state107_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state107_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state107_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state107_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state107_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state107_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state107_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state107_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state108_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state108_15_0 = reservoir_state[15] <<< 0;
wire signed [31:0] shifted_state108_15_1 = reservoir_state[15] <<< 1;
wire signed [31:0] shifted_state108_15_3 = reservoir_state[15] <<< 3;
wire signed [31:0] shifted_state108_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state108_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state108_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state108_19_1 = reservoir_state[19] <<< 1;
wire signed [31:0] shifted_state108_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state108_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state108_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state108_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state108_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state108_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state108_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state108_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state108_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state108_39_0 = reservoir_state[39] <<< 0;
wire signed [31:0] shifted_state108_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state108_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state108_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state108_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state108_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state108_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state108_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state108_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state108_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state108_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state108_67_2 = reservoir_state[67] <<< 2;
wire signed [31:0] shifted_state108_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state108_67_6 = reservoir_state[67] <<< 6;
wire signed [31:0] shifted_state108_67_7 = reservoir_state[67] <<< 7;
wire signed [31:0] shifted_state108_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state108_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state108_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state108_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state108_91_1 = reservoir_state[91] <<< 1;
wire signed [31:0] shifted_state108_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state108_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state108_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state108_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state108_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state108_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state108_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state108_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state108_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state108_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state108_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state108_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state108_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state108_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state108_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state108_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state108_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state108_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state108_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state108_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state108_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state108_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state108_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state108_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state108_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state108_151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state108_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state108_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state108_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state108_159_1 = reservoir_state[159] <<< 1;
wire signed [31:0] shifted_state108_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state108_159_5 = reservoir_state[159] <<< 5;
wire signed [31:0] shifted_state108_159_6 = reservoir_state[159] <<< 6;
wire signed [31:0] shifted_state108_159_7 = reservoir_state[159] <<< 7;
wire signed [31:0] shifted_state108_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state108_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state108_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state108_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state108_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state108_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state108_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state108_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state108_182_1 = reservoir_state[182] <<< 1;
wire signed [31:0] shifted_state108_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state108_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state108_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state108_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state108_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state108_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state109_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state109_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state109_1_3 = reservoir_state[1] <<< 3;
wire signed [31:0] shifted_state109_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state109_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state109_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state109_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state109_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state109_13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state109_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state109_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state109_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state109_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state109_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state109_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state109_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state109_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state109_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state109_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state109_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state109_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state109_55_2 = reservoir_state[55] <<< 2;
wire signed [31:0] shifted_state109_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state109_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state109_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state109_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state109_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state109_90_4 = reservoir_state[90] <<< 4;
wire signed [31:0] shifted_state109_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state109_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state109_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state109_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state109_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state109_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state109_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state109_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state109_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state109_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state109_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state109_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state109_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state109_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state109_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state109_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state109_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state109_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state109_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state109_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state109_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state109_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state109_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state109_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state109_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state109_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state109_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state109_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state109_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state109_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state109_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state109_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state109_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state109_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state109_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state109_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state109_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state109_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state109_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state109_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state109_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state109_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state109_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state109_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state109_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state109_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state110_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state110_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state110_15_0 = reservoir_state[15] <<< 0;
wire signed [31:0] shifted_state110_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state110_15_3 = reservoir_state[15] <<< 3;
wire signed [31:0] shifted_state110_15_4 = reservoir_state[15] <<< 4;
wire signed [31:0] shifted_state110_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state110_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state110_30_5 = reservoir_state[30] <<< 5;
wire signed [31:0] shifted_state110_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state110_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state110_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state110_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state110_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state110_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state110_58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state110_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state110_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state110_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state110_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state110_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state110_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state110_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state110_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state110_65_4 = reservoir_state[65] <<< 4;
wire signed [31:0] shifted_state110_68_1 = reservoir_state[68] <<< 1;
wire signed [31:0] shifted_state110_68_2 = reservoir_state[68] <<< 2;
wire signed [31:0] shifted_state110_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state110_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state110_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state110_70_4 = reservoir_state[70] <<< 4;
wire signed [31:0] shifted_state110_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state110_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state110_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state110_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state110_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state110_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state110_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state110_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state110_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state110_85_3 = reservoir_state[85] <<< 3;
wire signed [31:0] shifted_state110_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state110_114_2 = reservoir_state[114] <<< 2;
wire signed [31:0] shifted_state110_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state110_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state110_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state110_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state110_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state110_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state110_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state110_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state110_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state110_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state110_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state110_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state110_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state110_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state110_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state110_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state110_147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state110_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state110_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state110_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state110_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state110_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state110_161_0 = reservoir_state[161] <<< 0;
wire signed [31:0] shifted_state110_161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state110_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state110_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state110_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state110_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state110_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state110_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state110_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state110_171_6 = reservoir_state[171] <<< 6;
wire signed [31:0] shifted_state110_171_7 = reservoir_state[171] <<< 7;
wire signed [31:0] shifted_state110_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state110_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state110_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state110_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state110_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state110_179_2 = reservoir_state[179] <<< 2;
wire signed [31:0] shifted_state110_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state110_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state110_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state110_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state110_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state110_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state110_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state110_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state110_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state110_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state110_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state110_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state110_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state110_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state110_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state110_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state111_15_1 = reservoir_state[15] <<< 1;
wire signed [31:0] shifted_state111_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state111_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state111_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state111_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state111_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state111_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state111_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state111_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state111_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state111_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state111_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state111_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state111_84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state111_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state111_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state111_90_4 = reservoir_state[90] <<< 4;
wire signed [31:0] shifted_state111_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state111_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state111_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state111_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state111_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state111_93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state111_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state111_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state111_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state111_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state111_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state111_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state111_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state111_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state111_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state111_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state111_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state111_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state111_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state111_134_2 = reservoir_state[134] <<< 2;
wire signed [31:0] shifted_state111_134_4 = reservoir_state[134] <<< 4;
wire signed [31:0] shifted_state111_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state111_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state111_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state111_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state111_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state111_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state111_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state111_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state111_169_2 = reservoir_state[169] <<< 2;
wire signed [31:0] shifted_state111_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state111_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state111_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state111_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state111_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state111_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state111_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state111_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state111_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state111_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state111_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state112_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state112_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state112_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state112_34_2 = reservoir_state[34] <<< 2;
wire signed [31:0] shifted_state112_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state112_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state112_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state112_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state112_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state112_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state112_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state112_65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state112_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state112_65_5 = reservoir_state[65] <<< 5;
wire signed [31:0] shifted_state112_65_6 = reservoir_state[65] <<< 6;
wire signed [31:0] shifted_state112_65_7 = reservoir_state[65] <<< 7;
wire signed [31:0] shifted_state112_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state112_68_1 = reservoir_state[68] <<< 1;
wire signed [31:0] shifted_state112_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state112_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state112_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state112_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state112_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state112_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state112_92_1 = reservoir_state[92] <<< 1;
wire signed [31:0] shifted_state112_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state112_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state112_92_4 = reservoir_state[92] <<< 4;
wire signed [31:0] shifted_state112_119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state112_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state112_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state112_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state112_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state112_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state112_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state112_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state112_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state112_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state112_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state112_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state112_135_4 = reservoir_state[135] <<< 4;
wire signed [31:0] shifted_state112_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state112_135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state112_135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state112_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state112_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state112_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state112_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state112_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state112_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state112_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state112_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state112_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state112_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state112_173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state112_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state112_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state112_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state112_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state112_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state112_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state112_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state113_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state113_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state113_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state113_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state113_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state113_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state113_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state113_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state113_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state113_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state113_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state113_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state113_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state113_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state113_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state113_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state113_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state113_40_5 = reservoir_state[40] <<< 5;
wire signed [31:0] shifted_state113_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state113_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state113_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state113_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state113_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state113_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state113_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state113_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state113_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state113_84_2 = reservoir_state[84] <<< 2;
wire signed [31:0] shifted_state113_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state113_84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state113_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state113_87_3 = reservoir_state[87] <<< 3;
wire signed [31:0] shifted_state113_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state113_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state113_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state113_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state113_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state113_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state113_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state113_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state113_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state113_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state113_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state113_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state113_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state113_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state113_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state113_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state113_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state113_136_2 = reservoir_state[136] <<< 2;
wire signed [31:0] shifted_state113_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state113_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state113_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state113_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state113_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state113_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state113_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state113_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state113_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state113_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state113_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state113_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state113_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state113_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state113_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state113_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state113_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state113_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state113_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state113_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state113_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state113_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state113_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state113_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state113_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state114_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state114_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state114_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state114_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state114_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state114_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state114_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state114_5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state114_5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state114_5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state114_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state114_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state114_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state114_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state114_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state114_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state114_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state114_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state114_29_1 = reservoir_state[29] <<< 1;
wire signed [31:0] shifted_state114_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state114_29_5 = reservoir_state[29] <<< 5;
wire signed [31:0] shifted_state114_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state114_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state114_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state114_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state114_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state114_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state114_39_0 = reservoir_state[39] <<< 0;
wire signed [31:0] shifted_state114_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state114_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state114_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state114_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state114_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state114_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state114_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state114_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state114_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state114_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state114_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state114_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state114_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state114_58_2 = reservoir_state[58] <<< 2;
wire signed [31:0] shifted_state114_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state114_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state114_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state114_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state114_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state114_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state114_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state114_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state114_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state114_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state114_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state114_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state114_108_4 = reservoir_state[108] <<< 4;
wire signed [31:0] shifted_state114_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state114_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state114_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state114_110_2 = reservoir_state[110] <<< 2;
wire signed [31:0] shifted_state114_110_3 = reservoir_state[110] <<< 3;
wire signed [31:0] shifted_state114_110_4 = reservoir_state[110] <<< 4;
wire signed [31:0] shifted_state114_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state114_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state114_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state114_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state114_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state114_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state114_126_3 = reservoir_state[126] <<< 3;
wire signed [31:0] shifted_state114_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state114_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state114_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state114_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state114_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state114_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state114_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state114_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state114_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state115_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state115_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state115_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state115_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state115_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state115_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state115_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state115_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state115_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state115_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state115_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state115_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state115_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state115_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state115_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state115_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state115_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state115_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state115_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state115_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state115_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state115_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state115_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state115_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state115_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state115_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state115_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state115_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state115_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state115_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state115_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state115_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state115_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state115_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state115_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state115_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state115_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state115_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state115_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state115_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state115_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state115_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state115_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state115_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state115_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state115_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state115_88_5 = reservoir_state[88] <<< 5;
wire signed [31:0] shifted_state115_88_6 = reservoir_state[88] <<< 6;
wire signed [31:0] shifted_state115_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state115_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state115_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state115_101_2 = reservoir_state[101] <<< 2;
wire signed [31:0] shifted_state115_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state115_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state115_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state115_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state115_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state115_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state115_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state115_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state115_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state115_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state115_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state115_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state115_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state115_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state115_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state115_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state115_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state115_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state115_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state115_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state115_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state115_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state115_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state115_176_0 = reservoir_state[176] <<< 0;
wire signed [31:0] shifted_state115_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state115_176_2 = reservoir_state[176] <<< 2;
wire signed [31:0] shifted_state115_176_4 = reservoir_state[176] <<< 4;
wire signed [31:0] shifted_state115_176_5 = reservoir_state[176] <<< 5;
wire signed [31:0] shifted_state115_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state115_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state115_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state115_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state115_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state115_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state115_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state115_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state115_185_0 = reservoir_state[185] <<< 0;
wire signed [31:0] shifted_state115_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state115_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state115_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state115_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state115_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state115_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state115_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state115_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state115_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state115_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state115_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state116_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state116_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state116_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state116_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state116_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state116_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state116_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state116_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state116_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state116_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state116_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state116_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state116_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state116_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state116_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state116_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state116_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state116_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state116_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state116_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state116_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state116_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state116_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state116_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state116_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state116_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state116_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state116_29_2 = reservoir_state[29] <<< 2;
wire signed [31:0] shifted_state116_29_3 = reservoir_state[29] <<< 3;
wire signed [31:0] shifted_state116_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state116_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state116_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state116_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state116_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state116_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state116_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state116_73_3 = reservoir_state[73] <<< 3;
wire signed [31:0] shifted_state116_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state116_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state116_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state116_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state116_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state116_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state116_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state116_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state116_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state116_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state116_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state116_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state116_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state116_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state116_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state116_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state116_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state116_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state116_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state116_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state116_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state116_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state116_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state116_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state116_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state116_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state116_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state116_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state116_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state116_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state116_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state116_154_0 = reservoir_state[154] <<< 0;
wire signed [31:0] shifted_state116_154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state116_154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state116_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state116_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state116_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state116_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state116_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state116_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state116_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state116_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state116_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state116_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state116_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state116_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state116_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state116_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state116_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state116_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state116_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state116_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state116_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state117_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state117_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state117_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state117_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state117_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state117_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state117_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state117_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state117_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state117_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state117_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state117_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state117_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state117_36_4 = reservoir_state[36] <<< 4;
wire signed [31:0] shifted_state117_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state117_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state117_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state117_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state117_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state117_68_2 = reservoir_state[68] <<< 2;
wire signed [31:0] shifted_state117_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state117_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state117_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state117_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state117_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state117_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state117_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state117_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state117_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state117_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state117_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state117_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state117_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state117_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state117_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state117_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state117_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state117_101_2 = reservoir_state[101] <<< 2;
wire signed [31:0] shifted_state117_101_3 = reservoir_state[101] <<< 3;
wire signed [31:0] shifted_state117_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state117_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state117_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state117_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state117_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state117_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state117_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state117_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state117_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state117_144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state117_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state117_144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state117_144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state117_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state117_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state117_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state117_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state117_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state117_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state117_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state117_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state117_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state117_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state117_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state117_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state117_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state117_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state117_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state118_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state118_1_3 = reservoir_state[1] <<< 3;
wire signed [31:0] shifted_state118_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state118_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state118_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state118_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state118_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state118_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state118_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state118_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state118_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state118_9_0 = reservoir_state[9] <<< 0;
wire signed [31:0] shifted_state118_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state118_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state118_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state118_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state118_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state118_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state118_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state118_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state118_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state118_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state118_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state118_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state118_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state118_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state118_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state118_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state118_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state118_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state118_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state118_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state118_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state118_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state118_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state118_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state118_65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state118_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state118_65_2 = reservoir_state[65] <<< 2;
wire signed [31:0] shifted_state118_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state118_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state118_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state118_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state118_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state118_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state118_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state118_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state118_85_7 = reservoir_state[85] <<< 7;
wire signed [31:0] shifted_state118_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state118_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state118_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state118_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state118_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state118_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state118_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state118_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state118_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state118_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state118_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state118_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state118_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state118_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state118_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state118_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state118_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state118_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state118_147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state118_147_5 = reservoir_state[147] <<< 5;
wire signed [31:0] shifted_state118_147_6 = reservoir_state[147] <<< 6;
wire signed [31:0] shifted_state118_147_7 = reservoir_state[147] <<< 7;
wire signed [31:0] shifted_state118_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state118_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state118_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state118_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state119_3_1 = reservoir_state[3] <<< 1;
wire signed [31:0] shifted_state119_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state119_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state119_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state119_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state119_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state119_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state119_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state119_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state119_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state119_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state119_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state119_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state119_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state119_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state119_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state119_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state119_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state119_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state119_51_6 = reservoir_state[51] <<< 6;
wire signed [31:0] shifted_state119_51_7 = reservoir_state[51] <<< 7;
wire signed [31:0] shifted_state119_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state119_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state119_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state119_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state119_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state119_56_2 = reservoir_state[56] <<< 2;
wire signed [31:0] shifted_state119_56_5 = reservoir_state[56] <<< 5;
wire signed [31:0] shifted_state119_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state119_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state119_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state119_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state119_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state119_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state119_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state119_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state119_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state119_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state119_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state119_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state119_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state119_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state119_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state119_103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state119_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state119_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state119_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state119_124_6 = reservoir_state[124] <<< 6;
wire signed [31:0] shifted_state119_124_7 = reservoir_state[124] <<< 7;
wire signed [31:0] shifted_state119_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state119_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state119_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state119_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state119_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state119_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state119_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state119_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state119_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state119_167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state119_167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state119_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state119_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state119_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state119_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state119_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state119_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state119_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state119_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state119_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state119_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state119_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state119_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state120_2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state120_2_3 = reservoir_state[2] <<< 3;
wire signed [31:0] shifted_state120_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state120_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state120_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state120_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state120_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state120_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state120_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state120_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state120_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state120_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state120_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state120_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state120_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state120_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state120_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state120_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state120_48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state120_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state120_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state120_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state120_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state120_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state120_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state120_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state120_70_2 = reservoir_state[70] <<< 2;
wire signed [31:0] shifted_state120_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state120_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state120_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state120_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state120_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state120_74_3 = reservoir_state[74] <<< 3;
wire signed [31:0] shifted_state120_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state120_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state120_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state120_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state120_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state120_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state120_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state120_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state120_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state120_98_5 = reservoir_state[98] <<< 5;
wire signed [31:0] shifted_state120_98_6 = reservoir_state[98] <<< 6;
wire signed [31:0] shifted_state120_98_7 = reservoir_state[98] <<< 7;
wire signed [31:0] shifted_state120_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state120_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state120_124_2 = reservoir_state[124] <<< 2;
wire signed [31:0] shifted_state120_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state120_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state120_124_6 = reservoir_state[124] <<< 6;
wire signed [31:0] shifted_state120_124_7 = reservoir_state[124] <<< 7;
wire signed [31:0] shifted_state120_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state120_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state120_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state120_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state120_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state120_171_0 = reservoir_state[171] <<< 0;
wire signed [31:0] shifted_state120_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state120_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state120_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state120_171_5 = reservoir_state[171] <<< 5;
wire signed [31:0] shifted_state120_171_6 = reservoir_state[171] <<< 6;
wire signed [31:0] shifted_state120_171_7 = reservoir_state[171] <<< 7;
wire signed [31:0] shifted_state120_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state120_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state120_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state120_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state120_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state120_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state120_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state120_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state120_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state120_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state120_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state121_14_0 = reservoir_state[14] <<< 0;
wire signed [31:0] shifted_state121_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state121_14_3 = reservoir_state[14] <<< 3;
wire signed [31:0] shifted_state121_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state121_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state121_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state121_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state121_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state121_70_0 = reservoir_state[70] <<< 0;
wire signed [31:0] shifted_state121_70_2 = reservoir_state[70] <<< 2;
wire signed [31:0] shifted_state121_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state121_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state121_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state121_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state121_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state121_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state121_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state121_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state121_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state121_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state121_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state121_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state121_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state121_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state121_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state121_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state121_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state121_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state121_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state121_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state121_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state121_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state121_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state121_185_0 = reservoir_state[185] <<< 0;
wire signed [31:0] shifted_state121_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state121_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state121_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state121_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state121_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state121_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state121_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state121_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state121_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state121_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state122_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state122_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state122_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state122_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state122_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state122_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state122_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state122_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state122_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state122_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state122_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state122_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state122_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state122_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state122_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state122_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state122_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state122_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state122_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state122_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state122_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state122_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state122_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state122_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state122_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state122_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state122_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state122_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state122_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state122_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state122_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state122_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state122_55_2 = reservoir_state[55] <<< 2;
wire signed [31:0] shifted_state122_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state122_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state122_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state122_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state122_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state122_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state122_91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state122_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state122_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state122_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state122_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state122_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state122_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state122_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state122_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state122_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state122_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state122_112_3 = reservoir_state[112] <<< 3;
wire signed [31:0] shifted_state122_114_2 = reservoir_state[114] <<< 2;
wire signed [31:0] shifted_state122_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state122_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state122_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state122_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state122_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state122_143_0 = reservoir_state[143] <<< 0;
wire signed [31:0] shifted_state122_143_3 = reservoir_state[143] <<< 3;
wire signed [31:0] shifted_state122_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state122_143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state122_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state122_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state122_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state122_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state122_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state122_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state122_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state122_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state122_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state122_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state122_182_1 = reservoir_state[182] <<< 1;
wire signed [31:0] shifted_state122_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state122_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state122_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state122_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state122_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state122_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state122_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state122_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state122_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state122_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state122_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state122_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state122_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state122_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state122_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state122_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state122_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state122_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state122_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state122_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state122_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state123_2_0 = reservoir_state[2] <<< 0;
wire signed [31:0] shifted_state123_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state123_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state123_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state123_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state123_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state123_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state123_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state123_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state123_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state123_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state123_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state123_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state123_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state123_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state123_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state123_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state123_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state123_48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state123_48_6 = reservoir_state[48] <<< 6;
wire signed [31:0] shifted_state123_48_7 = reservoir_state[48] <<< 7;
wire signed [31:0] shifted_state123_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state123_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state123_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state123_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state123_60_4 = reservoir_state[60] <<< 4;
wire signed [31:0] shifted_state123_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state123_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state123_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state123_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state123_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state123_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state123_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state123_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state123_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state123_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state123_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state123_72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state123_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state123_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state123_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state123_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state123_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state123_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state123_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state123_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state123_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state123_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state123_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state123_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state123_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state123_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state123_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state123_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state123_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state123_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state123_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state123_135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state123_135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state123_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state123_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state123_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state123_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state123_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state123_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state123_152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state123_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state123_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state123_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state123_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state123_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state123_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state123_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state123_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state123_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state123_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state123_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state123_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state123_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state123_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state124_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state124_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state124_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state124_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state124_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state124_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state124_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state124_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state124_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state124_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state124_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state124_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state124_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state124_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state124_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state124_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state124_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state124_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state124_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state124_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state124_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state124_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state124_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state124_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state124_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state124_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state124_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state124_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state124_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state124_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state124_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state124_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state124_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state124_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state124_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state124_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state124_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state124_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state124_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state124_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state124_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state124_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state124_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state124_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state124_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state124_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state124_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state124_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state124_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state124_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state124_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state124_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state124_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state124_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state124_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state124_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state124_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state124_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state124_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state124_119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state124_119_2 = reservoir_state[119] <<< 2;
wire signed [31:0] shifted_state124_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state124_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state124_119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state124_119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state124_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state124_136_2 = reservoir_state[136] <<< 2;
wire signed [31:0] shifted_state124_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state124_142_0 = reservoir_state[142] <<< 0;
wire signed [31:0] shifted_state124_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state124_142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state124_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state124_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state124_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state124_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state124_151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state124_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state124_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state124_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state124_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state124_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state124_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state124_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state124_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state124_162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state124_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state124_185_2 = reservoir_state[185] <<< 2;
wire signed [31:0] shifted_state124_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state124_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state124_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state124_186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state124_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state124_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state124_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state124_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state124_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state124_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state124_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state124_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state124_189_6 = reservoir_state[189] <<< 6;
wire signed [31:0] shifted_state124_189_7 = reservoir_state[189] <<< 7;
wire signed [31:0] shifted_state124_196_0 = reservoir_state[196] <<< 0;
wire signed [31:0] shifted_state124_196_3 = reservoir_state[196] <<< 3;
wire signed [31:0] shifted_state124_196_4 = reservoir_state[196] <<< 4;
wire signed [31:0] shifted_state124_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state124_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state125_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state125_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state125_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state125_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state125_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state125_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state125_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state125_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state125_8_6 = reservoir_state[8] <<< 6;
wire signed [31:0] shifted_state125_8_7 = reservoir_state[8] <<< 7;
wire signed [31:0] shifted_state125_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state125_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state125_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state125_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state125_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state125_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state125_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state125_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state125_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state125_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state125_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state125_64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state125_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state125_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state125_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state125_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state125_79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state125_79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state125_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state125_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state125_84_2 = reservoir_state[84] <<< 2;
wire signed [31:0] shifted_state125_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state125_84_5 = reservoir_state[84] <<< 5;
wire signed [31:0] shifted_state125_84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state125_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state125_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state125_90_4 = reservoir_state[90] <<< 4;
wire signed [31:0] shifted_state125_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state125_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state125_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state125_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state125_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state125_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state125_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state125_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state125_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state125_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state125_124_2 = reservoir_state[124] <<< 2;
wire signed [31:0] shifted_state125_124_3 = reservoir_state[124] <<< 3;
wire signed [31:0] shifted_state125_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state125_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state125_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state125_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state125_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state125_137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state125_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state125_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state125_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state125_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state125_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state125_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state125_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state125_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state125_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state125_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state125_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state125_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state125_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state125_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state125_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state125_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state125_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state125_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state125_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state125_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state126_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state126_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state126_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state126_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state126_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state126_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state126_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state126_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state126_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state126_40_2 = reservoir_state[40] <<< 2;
wire signed [31:0] shifted_state126_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state126_40_5 = reservoir_state[40] <<< 5;
wire signed [31:0] shifted_state126_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state126_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state126_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state126_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state126_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state126_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state126_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state126_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state126_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state126_81_2 = reservoir_state[81] <<< 2;
wire signed [31:0] shifted_state126_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state126_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state126_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state126_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state126_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state126_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state126_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state126_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state126_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state126_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state126_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state126_110_1 = reservoir_state[110] <<< 1;
wire signed [31:0] shifted_state126_110_2 = reservoir_state[110] <<< 2;
wire signed [31:0] shifted_state126_110_4 = reservoir_state[110] <<< 4;
wire signed [31:0] shifted_state126_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state126_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state126_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state126_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state126_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state126_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state126_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state126_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state126_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state126_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state126_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state126_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state126_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state126_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state126_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state126_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state126_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state126_151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state126_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state126_158_3 = reservoir_state[158] <<< 3;
wire signed [31:0] shifted_state126_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state126_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state126_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state126_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state126_160_4 = reservoir_state[160] <<< 4;
wire signed [31:0] shifted_state126_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state126_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state126_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state126_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state126_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state126_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state126_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state126_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state126_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state126_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state126_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state127_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state127_8_1 = reservoir_state[8] <<< 1;
wire signed [31:0] shifted_state127_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state127_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state127_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state127_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state127_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state127_17_4 = reservoir_state[17] <<< 4;
wire signed [31:0] shifted_state127_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state127_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state127_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state127_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state127_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state127_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state127_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state127_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state127_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state127_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state127_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state127_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state127_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state127_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state127_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state127_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state127_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state127_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state127_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state127_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state127_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state127_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state127_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state127_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state127_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state127_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state127_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state127_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state127_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state127_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state127_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state127_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state127_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state128_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state128_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state128_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state128_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state128_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state128_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state128_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state128_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state128_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state128_91_1 = reservoir_state[91] <<< 1;
wire signed [31:0] shifted_state128_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state128_91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state128_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state128_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state128_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state128_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state128_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state128_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state128_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state128_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state128_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state128_114_1 = reservoir_state[114] <<< 1;
wire signed [31:0] shifted_state128_114_2 = reservoir_state[114] <<< 2;
wire signed [31:0] shifted_state128_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state128_119_3 = reservoir_state[119] <<< 3;
wire signed [31:0] shifted_state128_128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state128_128_2 = reservoir_state[128] <<< 2;
wire signed [31:0] shifted_state128_128_3 = reservoir_state[128] <<< 3;
wire signed [31:0] shifted_state128_128_4 = reservoir_state[128] <<< 4;
wire signed [31:0] shifted_state128_128_5 = reservoir_state[128] <<< 5;
wire signed [31:0] shifted_state128_128_6 = reservoir_state[128] <<< 6;
wire signed [31:0] shifted_state128_128_7 = reservoir_state[128] <<< 7;
wire signed [31:0] shifted_state128_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state128_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state128_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state128_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state128_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state128_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state128_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state128_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state128_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state128_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state128_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state128_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state128_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state128_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state128_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state128_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state128_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state128_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state128_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state128_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state128_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state129_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state129_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state129_34_0 = reservoir_state[34] <<< 0;
wire signed [31:0] shifted_state129_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state129_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state129_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state129_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state129_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state129_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state129_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state129_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state129_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state129_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state129_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state129_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state129_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state129_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state129_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state129_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state129_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state129_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state129_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state129_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state129_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state129_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state129_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state129_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state129_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state129_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state129_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state129_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state129_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state129_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state129_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state129_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state129_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state129_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state129_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state129_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state129_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state129_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state129_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state129_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state129_153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state129_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state129_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state129_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state129_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state129_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state129_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state129_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state129_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state129_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state129_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state129_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state129_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state129_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state129_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state129_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state129_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state129_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state129_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state129_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state129_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state129_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state130_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state130_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state130_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state130_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state130_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state130_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state130_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state130_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state130_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state130_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state130_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state130_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state130_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state130_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state130_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state130_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state130_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state130_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state130_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state130_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state130_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state130_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state130_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state130_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state130_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state130_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state130_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state130_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state130_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state130_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state130_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state130_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state130_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state130_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state130_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state130_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state130_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state130_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state130_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state130_85_3 = reservoir_state[85] <<< 3;
wire signed [31:0] shifted_state130_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state130_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state130_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state130_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state130_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state130_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state130_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state130_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state130_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state130_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state130_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state130_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state130_118_3 = reservoir_state[118] <<< 3;
wire signed [31:0] shifted_state130_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state130_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state130_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state130_146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state130_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state130_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state130_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state130_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state130_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state130_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state130_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state130_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state130_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state130_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state130_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state130_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state130_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state130_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state130_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state130_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state130_181_1 = reservoir_state[181] <<< 1;
wire signed [31:0] shifted_state130_181_3 = reservoir_state[181] <<< 3;
wire signed [31:0] shifted_state130_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state130_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state130_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state130_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state130_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state130_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state130_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state130_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state130_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state130_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state130_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state130_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state131_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state131_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state131_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state131_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state131_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state131_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state131_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state131_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state131_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state131_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state131_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state131_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state131_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state131_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state131_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state131_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state131_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state131_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state131_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state131_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state131_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state131_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state131_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state131_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state131_56_5 = reservoir_state[56] <<< 5;
wire signed [31:0] shifted_state131_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state131_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state131_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state131_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state131_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state131_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state131_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state131_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state131_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state131_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state131_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state131_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state131_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state131_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state131_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state131_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state131_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state131_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state131_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state131_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state131_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state131_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state131_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state131_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state131_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state131_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state131_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state131_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state131_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state131_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state131_118_3 = reservoir_state[118] <<< 3;
wire signed [31:0] shifted_state131_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state131_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state131_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state131_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state131_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state131_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state131_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state131_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state131_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state131_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state131_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state131_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state131_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state131_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state131_134_2 = reservoir_state[134] <<< 2;
wire signed [31:0] shifted_state131_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state131_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state131_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state131_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state131_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state131_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state131_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state131_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state131_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state131_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state132_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state132_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state132_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state132_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state132_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state132_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state132_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state132_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state132_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state132_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state132_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state132_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state132_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state132_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state132_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state132_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state132_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state132_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state132_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state132_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state132_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state132_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state132_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state132_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state132_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state132_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state132_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state132_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state132_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state132_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state132_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state132_48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state132_48_6 = reservoir_state[48] <<< 6;
wire signed [31:0] shifted_state132_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state132_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state132_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state132_60_4 = reservoir_state[60] <<< 4;
wire signed [31:0] shifted_state132_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state132_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state132_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state132_65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state132_65_5 = reservoir_state[65] <<< 5;
wire signed [31:0] shifted_state132_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state132_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state132_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state132_102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state132_102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state132_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state132_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state132_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state132_126_3 = reservoir_state[126] <<< 3;
wire signed [31:0] shifted_state132_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state132_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state132_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state132_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state132_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state132_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state132_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state132_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state132_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state132_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state132_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state132_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state132_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state132_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state133_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state133_5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state133_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state133_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state133_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state133_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state133_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state133_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state133_40_2 = reservoir_state[40] <<< 2;
wire signed [31:0] shifted_state133_40_5 = reservoir_state[40] <<< 5;
wire signed [31:0] shifted_state133_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state133_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state133_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state133_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state133_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state133_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state133_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state133_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state133_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state133_68_1 = reservoir_state[68] <<< 1;
wire signed [31:0] shifted_state133_68_2 = reservoir_state[68] <<< 2;
wire signed [31:0] shifted_state133_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state133_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state133_68_6 = reservoir_state[68] <<< 6;
wire signed [31:0] shifted_state133_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state133_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state133_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state133_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state133_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state133_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state133_84_2 = reservoir_state[84] <<< 2;
wire signed [31:0] shifted_state133_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state133_84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state133_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state133_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state133_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state133_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state133_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state133_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state133_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state133_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state133_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state133_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state133_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state133_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state133_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state133_111_4 = reservoir_state[111] <<< 4;
wire signed [31:0] shifted_state133_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state133_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state133_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state133_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state133_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state133_156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state133_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state133_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state133_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state133_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state133_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state133_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state133_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state133_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state133_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state133_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state133_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state133_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state133_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state133_176_3 = reservoir_state[176] <<< 3;
wire signed [31:0] shifted_state133_176_5 = reservoir_state[176] <<< 5;
wire signed [31:0] shifted_state133_176_6 = reservoir_state[176] <<< 6;
wire signed [31:0] shifted_state133_176_7 = reservoir_state[176] <<< 7;
wire signed [31:0] shifted_state133_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state133_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state133_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state133_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state133_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state133_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state133_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state133_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state133_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state133_199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state133_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state133_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state134_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state134_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state134_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state134_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state134_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state134_15_1 = reservoir_state[15] <<< 1;
wire signed [31:0] shifted_state134_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state134_15_4 = reservoir_state[15] <<< 4;
wire signed [31:0] shifted_state134_15_5 = reservoir_state[15] <<< 5;
wire signed [31:0] shifted_state134_15_6 = reservoir_state[15] <<< 6;
wire signed [31:0] shifted_state134_15_7 = reservoir_state[15] <<< 7;
wire signed [31:0] shifted_state134_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state134_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state134_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state134_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state134_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state134_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state134_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state134_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state134_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state134_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state134_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state134_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state134_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state134_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state134_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state134_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state134_70_4 = reservoir_state[70] <<< 4;
wire signed [31:0] shifted_state134_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state134_88_5 = reservoir_state[88] <<< 5;
wire signed [31:0] shifted_state134_88_6 = reservoir_state[88] <<< 6;
wire signed [31:0] shifted_state134_88_7 = reservoir_state[88] <<< 7;
wire signed [31:0] shifted_state134_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state134_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state134_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state134_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state134_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state134_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state134_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state134_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state134_94_2 = reservoir_state[94] <<< 2;
wire signed [31:0] shifted_state134_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state134_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state134_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state134_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state134_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state134_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state134_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state134_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state134_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state134_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state134_108_1 = reservoir_state[108] <<< 1;
wire signed [31:0] shifted_state134_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state134_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state134_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state134_134_2 = reservoir_state[134] <<< 2;
wire signed [31:0] shifted_state134_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state134_134_5 = reservoir_state[134] <<< 5;
wire signed [31:0] shifted_state134_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state134_134_7 = reservoir_state[134] <<< 7;
wire signed [31:0] shifted_state134_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state134_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state134_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state134_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state134_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state134_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state134_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state134_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state134_194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state134_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state135_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state135_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state135_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state135_23_4 = reservoir_state[23] <<< 4;
wire signed [31:0] shifted_state135_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state135_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state135_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state135_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state135_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state135_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state135_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state135_65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state135_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state135_65_2 = reservoir_state[65] <<< 2;
wire signed [31:0] shifted_state135_65_3 = reservoir_state[65] <<< 3;
wire signed [31:0] shifted_state135_65_4 = reservoir_state[65] <<< 4;
wire signed [31:0] shifted_state135_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state135_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state135_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state135_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state135_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state135_81_2 = reservoir_state[81] <<< 2;
wire signed [31:0] shifted_state135_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state135_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state135_91_1 = reservoir_state[91] <<< 1;
wire signed [31:0] shifted_state135_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state135_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state135_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state135_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state135_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state135_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state135_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state135_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state135_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state135_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state135_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state135_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state135_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state135_142_0 = reservoir_state[142] <<< 0;
wire signed [31:0] shifted_state135_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state135_142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state135_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state135_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state135_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state135_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state135_144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state135_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state135_144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state135_144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state135_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state135_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state135_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state135_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state135_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state135_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state135_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state135_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state135_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state135_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state135_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state135_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state135_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state135_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state135_182_1 = reservoir_state[182] <<< 1;
wire signed [31:0] shifted_state135_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state135_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state135_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state135_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state135_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state135_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state135_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state135_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state135_191_3 = reservoir_state[191] <<< 3;
wire signed [31:0] shifted_state135_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state135_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state135_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state136_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state136_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state136_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state136_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state136_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state136_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state136_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state136_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state136_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state136_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state136_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state136_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state136_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state136_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state136_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state136_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state136_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state136_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state136_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state136_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state136_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state136_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state136_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state136_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state136_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state136_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state136_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state136_33_4 = reservoir_state[33] <<< 4;
wire signed [31:0] shifted_state136_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state136_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state136_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state136_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state136_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state136_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state136_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state136_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state136_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state136_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state136_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state136_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state136_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state136_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state136_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state136_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state136_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state136_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state136_53_1 = reservoir_state[53] <<< 1;
wire signed [31:0] shifted_state136_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state136_53_3 = reservoir_state[53] <<< 3;
wire signed [31:0] shifted_state136_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state136_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state136_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state136_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state136_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state136_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state136_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state136_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state136_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state136_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state136_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state136_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state136_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state136_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state136_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state136_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state136_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state136_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state136_85_7 = reservoir_state[85] <<< 7;
wire signed [31:0] shifted_state136_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state136_87_2 = reservoir_state[87] <<< 2;
wire signed [31:0] shifted_state136_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state136_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state136_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state136_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state136_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state136_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state136_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state136_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state136_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state136_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state136_120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state136_120_5 = reservoir_state[120] <<< 5;
wire signed [31:0] shifted_state136_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state136_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state136_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state136_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state136_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state136_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state136_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state136_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state136_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state136_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state136_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state136_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state136_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state136_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state136_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state136_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state136_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state136_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state136_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state136_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state136_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state136_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state136_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state136_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state136_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state137_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state137_8_5 = reservoir_state[8] <<< 5;
wire signed [31:0] shifted_state137_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state137_9_6 = reservoir_state[9] <<< 6;
wire signed [31:0] shifted_state137_9_7 = reservoir_state[9] <<< 7;
wire signed [31:0] shifted_state137_23_4 = reservoir_state[23] <<< 4;
wire signed [31:0] shifted_state137_23_5 = reservoir_state[23] <<< 5;
wire signed [31:0] shifted_state137_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state137_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state137_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state137_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state137_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state137_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state137_40_5 = reservoir_state[40] <<< 5;
wire signed [31:0] shifted_state137_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state137_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state137_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state137_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state137_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state137_51_6 = reservoir_state[51] <<< 6;
wire signed [31:0] shifted_state137_51_7 = reservoir_state[51] <<< 7;
wire signed [31:0] shifted_state137_52_1 = reservoir_state[52] <<< 1;
wire signed [31:0] shifted_state137_52_4 = reservoir_state[52] <<< 4;
wire signed [31:0] shifted_state137_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state137_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state137_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state137_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state137_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state137_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state137_66_2 = reservoir_state[66] <<< 2;
wire signed [31:0] shifted_state137_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state137_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state137_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state137_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state137_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state137_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state137_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state137_92_4 = reservoir_state[92] <<< 4;
wire signed [31:0] shifted_state137_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state137_92_6 = reservoir_state[92] <<< 6;
wire signed [31:0] shifted_state137_92_7 = reservoir_state[92] <<< 7;
wire signed [31:0] shifted_state137_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state137_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state137_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state137_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state137_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state137_103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state137_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state137_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state137_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state137_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state137_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state137_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state137_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state137_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state137_112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state137_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state137_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state137_114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state137_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state137_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state137_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state137_115_4 = reservoir_state[115] <<< 4;
wire signed [31:0] shifted_state137_115_6 = reservoir_state[115] <<< 6;
wire signed [31:0] shifted_state137_115_7 = reservoir_state[115] <<< 7;
wire signed [31:0] shifted_state137_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state137_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state137_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state137_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state137_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state137_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state137_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state137_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state137_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state137_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state137_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state137_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state137_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state137_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state137_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state137_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state137_182_1 = reservoir_state[182] <<< 1;
wire signed [31:0] shifted_state137_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state137_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state137_188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state137_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state137_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state137_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state137_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state137_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state137_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state138_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state138_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state138_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state138_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state138_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state138_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state138_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state138_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state138_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state138_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state138_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state138_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state138_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state138_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state138_72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state138_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state138_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state138_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state138_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state138_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state138_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state138_81_2 = reservoir_state[81] <<< 2;
wire signed [31:0] shifted_state138_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state138_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state138_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state138_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state138_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state138_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state138_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state138_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state138_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state138_85_7 = reservoir_state[85] <<< 7;
wire signed [31:0] shifted_state138_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state138_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state138_94_2 = reservoir_state[94] <<< 2;
wire signed [31:0] shifted_state138_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state138_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state138_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state138_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state138_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state138_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state138_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state138_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state138_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state138_125_4 = reservoir_state[125] <<< 4;
wire signed [31:0] shifted_state138_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state138_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state138_140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state138_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state138_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state138_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state138_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state138_144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state138_144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state138_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state138_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state138_149_5 = reservoir_state[149] <<< 5;
wire signed [31:0] shifted_state138_149_6 = reservoir_state[149] <<< 6;
wire signed [31:0] shifted_state138_149_7 = reservoir_state[149] <<< 7;
wire signed [31:0] shifted_state138_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state138_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state138_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state138_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state138_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state138_158_3 = reservoir_state[158] <<< 3;
wire signed [31:0] shifted_state138_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state138_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state138_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state138_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state138_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state138_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state138_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state138_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state138_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state138_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state138_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state138_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state138_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state138_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state138_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state138_183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state138_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state138_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state138_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state138_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state138_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state138_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state138_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state138_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state139_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state139_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state139_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state139_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state139_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state139_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state139_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state139_49_4 = reservoir_state[49] <<< 4;
wire signed [31:0] shifted_state139_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state139_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state139_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state139_56_0 = reservoir_state[56] <<< 0;
wire signed [31:0] shifted_state139_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state139_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state139_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state139_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state139_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state139_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state139_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state139_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state139_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state139_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state139_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state139_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state139_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state139_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state139_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state139_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state139_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state139_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state139_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state139_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state139_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state139_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state139_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state139_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state139_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state139_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state139_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state139_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state139_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state139_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state139_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state139_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state139_151_4 = reservoir_state[151] <<< 4;
wire signed [31:0] shifted_state139_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state139_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state139_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state139_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state139_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state139_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state139_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state139_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state139_185_0 = reservoir_state[185] <<< 0;
wire signed [31:0] shifted_state139_185_2 = reservoir_state[185] <<< 2;
wire signed [31:0] shifted_state139_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state139_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state139_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state140_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state140_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state140_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state140_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state140_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state140_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state140_27_4 = reservoir_state[27] <<< 4;
wire signed [31:0] shifted_state140_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state140_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state140_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state140_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state140_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state140_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state140_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state140_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state140_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state140_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state140_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state140_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state140_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state140_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state140_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state140_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state140_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state140_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state140_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state140_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state140_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state140_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state140_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state140_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state140_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state140_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state140_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state140_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state140_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state140_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state140_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state140_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state140_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state140_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state140_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state140_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state140_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state140_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state140_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state140_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state140_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state140_152_0 = reservoir_state[152] <<< 0;
wire signed [31:0] shifted_state140_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state140_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state140_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state140_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state140_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state140_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state140_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state140_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state140_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state140_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state140_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state140_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state140_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state140_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state140_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state140_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state140_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state140_182_1 = reservoir_state[182] <<< 1;
wire signed [31:0] shifted_state140_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state140_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state140_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state140_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state141_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state141_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state141_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state141_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state141_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state141_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state141_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state141_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state141_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state141_13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state141_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state141_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state141_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state141_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state141_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state141_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state141_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state141_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state141_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state141_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state141_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state141_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state141_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state141_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state141_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state141_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state141_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state141_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state141_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state141_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state141_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state141_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state141_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state141_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state141_65_6 = reservoir_state[65] <<< 6;
wire signed [31:0] shifted_state141_65_7 = reservoir_state[65] <<< 7;
wire signed [31:0] shifted_state141_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state141_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state141_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state141_85_3 = reservoir_state[85] <<< 3;
wire signed [31:0] shifted_state141_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state141_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state141_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state141_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state141_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state141_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state141_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state141_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state141_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state141_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state141_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state141_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state141_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state141_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state141_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state141_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state141_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state141_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state141_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state141_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state141_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state141_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state141_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state141_131_2 = reservoir_state[131] <<< 2;
wire signed [31:0] shifted_state141_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state141_131_5 = reservoir_state[131] <<< 5;
wire signed [31:0] shifted_state141_148_4 = reservoir_state[148] <<< 4;
wire signed [31:0] shifted_state141_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state141_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state141_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state141_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state141_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state141_151_0 = reservoir_state[151] <<< 0;
wire signed [31:0] shifted_state141_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state141_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state141_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state141_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state141_160_2 = reservoir_state[160] <<< 2;
wire signed [31:0] shifted_state141_160_4 = reservoir_state[160] <<< 4;
wire signed [31:0] shifted_state141_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state141_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state141_171_0 = reservoir_state[171] <<< 0;
wire signed [31:0] shifted_state141_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state141_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state141_171_6 = reservoir_state[171] <<< 6;
wire signed [31:0] shifted_state141_171_7 = reservoir_state[171] <<< 7;
wire signed [31:0] shifted_state141_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state141_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state141_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state141_184_4 = reservoir_state[184] <<< 4;
wire signed [31:0] shifted_state141_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state141_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state141_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state141_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state141_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state141_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state141_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state141_197_0 = reservoir_state[197] <<< 0;
wire signed [31:0] shifted_state141_197_5 = reservoir_state[197] <<< 5;
wire signed [31:0] shifted_state141_197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state141_197_7 = reservoir_state[197] <<< 7;
wire signed [31:0] shifted_state142_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state142_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state142_5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state142_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state142_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state142_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state142_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state142_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state142_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state142_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state142_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state142_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state142_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state142_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state142_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state142_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state142_49_3 = reservoir_state[49] <<< 3;
wire signed [31:0] shifted_state142_49_4 = reservoir_state[49] <<< 4;
wire signed [31:0] shifted_state142_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state142_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state142_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state142_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state142_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state142_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state142_53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state142_53_1 = reservoir_state[53] <<< 1;
wire signed [31:0] shifted_state142_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state142_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state142_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state142_65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state142_65_3 = reservoir_state[65] <<< 3;
wire signed [31:0] shifted_state142_65_4 = reservoir_state[65] <<< 4;
wire signed [31:0] shifted_state142_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state142_71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state142_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state142_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state142_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state142_73_1 = reservoir_state[73] <<< 1;
wire signed [31:0] shifted_state142_73_2 = reservoir_state[73] <<< 2;
wire signed [31:0] shifted_state142_73_3 = reservoir_state[73] <<< 3;
wire signed [31:0] shifted_state142_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state142_73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state142_73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state142_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state142_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state142_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state142_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state142_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state142_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state142_84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state142_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state142_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state142_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state142_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state142_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state142_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state142_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state142_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state142_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state142_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state142_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state142_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state142_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state142_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state142_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state142_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state142_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state142_125_4 = reservoir_state[125] <<< 4;
wire signed [31:0] shifted_state142_125_5 = reservoir_state[125] <<< 5;
wire signed [31:0] shifted_state142_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state142_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state142_131_4 = reservoir_state[131] <<< 4;
wire signed [31:0] shifted_state142_131_6 = reservoir_state[131] <<< 6;
wire signed [31:0] shifted_state142_131_7 = reservoir_state[131] <<< 7;
wire signed [31:0] shifted_state142_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state142_138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state142_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state142_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state142_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state142_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state142_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state142_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state142_156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state142_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state142_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state142_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state142_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state142_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state142_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state142_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state142_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state142_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state142_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state142_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state142_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state142_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state142_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state142_196_3 = reservoir_state[196] <<< 3;
wire signed [31:0] shifted_state142_196_5 = reservoir_state[196] <<< 5;
wire signed [31:0] shifted_state143_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state143_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state143_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state143_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state143_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state143_9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state143_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state143_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state143_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state143_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state143_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state143_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state143_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state143_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state143_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state143_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state143_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state143_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state143_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state143_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state143_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state143_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state143_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state143_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state143_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state143_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state143_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state143_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state143_33_4 = reservoir_state[33] <<< 4;
wire signed [31:0] shifted_state143_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state143_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state143_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state143_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state143_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state143_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state143_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state143_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state143_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state143_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state143_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state143_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state143_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state143_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state143_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state143_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state143_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state143_103_0 = reservoir_state[103] <<< 0;
wire signed [31:0] shifted_state143_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state143_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state143_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state143_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state143_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state143_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state143_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state143_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state143_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state143_113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state143_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state143_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state143_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state143_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state143_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state143_134_2 = reservoir_state[134] <<< 2;
wire signed [31:0] shifted_state143_134_5 = reservoir_state[134] <<< 5;
wire signed [31:0] shifted_state143_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state143_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state143_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state143_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state143_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state143_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state143_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state143_183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state143_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state143_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state143_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state143_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state143_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state143_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state144_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state144_14_3 = reservoir_state[14] <<< 3;
wire signed [31:0] shifted_state144_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state144_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state144_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state144_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state144_15_0 = reservoir_state[15] <<< 0;
wire signed [31:0] shifted_state144_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state144_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state144_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state144_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state144_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state144_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state144_49_1 = reservoir_state[49] <<< 1;
wire signed [31:0] shifted_state144_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state144_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state144_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state144_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state144_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state144_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state144_51_6 = reservoir_state[51] <<< 6;
wire signed [31:0] shifted_state144_51_7 = reservoir_state[51] <<< 7;
wire signed [31:0] shifted_state144_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state144_84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state144_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state144_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state144_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state144_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state144_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state144_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state144_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state144_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state144_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state144_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state144_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state144_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state144_125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state144_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state144_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state144_128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state144_128_2 = reservoir_state[128] <<< 2;
wire signed [31:0] shifted_state144_134_4 = reservoir_state[134] <<< 4;
wire signed [31:0] shifted_state144_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state144_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state144_135_2 = reservoir_state[135] <<< 2;
wire signed [31:0] shifted_state144_135_3 = reservoir_state[135] <<< 3;
wire signed [31:0] shifted_state144_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state144_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state144_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state144_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state144_142_0 = reservoir_state[142] <<< 0;
wire signed [31:0] shifted_state144_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state144_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state144_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state144_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state144_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state144_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state144_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state144_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state144_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state144_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state144_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state144_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state144_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state144_181_1 = reservoir_state[181] <<< 1;
wire signed [31:0] shifted_state144_181_3 = reservoir_state[181] <<< 3;
wire signed [31:0] shifted_state144_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state144_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state144_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state144_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state144_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state145_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state145_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state145_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state145_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state145_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state145_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state145_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state145_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state145_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state145_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state145_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state145_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state145_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state145_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state145_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state145_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state145_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state145_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state145_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state145_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state145_49_4 = reservoir_state[49] <<< 4;
wire signed [31:0] shifted_state145_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state145_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state145_68_1 = reservoir_state[68] <<< 1;
wire signed [31:0] shifted_state145_68_2 = reservoir_state[68] <<< 2;
wire signed [31:0] shifted_state145_68_4 = reservoir_state[68] <<< 4;
wire signed [31:0] shifted_state145_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state145_68_7 = reservoir_state[68] <<< 7;
wire signed [31:0] shifted_state145_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state145_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state145_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state145_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state145_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state145_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state145_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state145_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state145_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state145_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state145_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state145_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state145_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state145_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state145_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state145_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state145_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state145_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state145_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state145_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state145_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state145_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state145_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state145_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state145_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state145_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state145_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state145_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state145_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state145_167_0 = reservoir_state[167] <<< 0;
wire signed [31:0] shifted_state145_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state145_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state145_167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state145_181_0 = reservoir_state[181] <<< 0;
wire signed [31:0] shifted_state145_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state145_181_3 = reservoir_state[181] <<< 3;
wire signed [31:0] shifted_state145_181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state145_181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state145_181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state145_181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state145_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state145_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state145_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state145_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state145_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state145_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state145_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state145_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state145_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state145_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state145_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state145_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state145_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state145_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state145_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state145_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state145_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state145_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state145_199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state145_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state145_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state145_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state146_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state146_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state146_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state146_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state146_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state146_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state146_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state146_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state146_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state146_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state146_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state146_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state146_33_3 = reservoir_state[33] <<< 3;
wire signed [31:0] shifted_state146_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state146_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state146_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state146_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state146_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state146_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state146_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state146_49_4 = reservoir_state[49] <<< 4;
wire signed [31:0] shifted_state146_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state146_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state146_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state146_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state146_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state146_66_2 = reservoir_state[66] <<< 2;
wire signed [31:0] shifted_state146_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state146_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state146_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state146_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state146_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state146_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state146_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state146_84_2 = reservoir_state[84] <<< 2;
wire signed [31:0] shifted_state146_84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state146_84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state146_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state146_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state146_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state146_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state146_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state146_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state146_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state146_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state146_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state146_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state146_119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state146_119_2 = reservoir_state[119] <<< 2;
wire signed [31:0] shifted_state146_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state146_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state146_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state146_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state146_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state146_184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state146_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state146_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state146_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state146_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state146_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state146_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state146_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state146_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state146_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state147_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state147_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state147_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state147_29_3 = reservoir_state[29] <<< 3;
wire signed [31:0] shifted_state147_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state147_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state147_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state147_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state147_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state147_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state147_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state147_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state147_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state147_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state147_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state147_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state147_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state147_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state147_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state147_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state147_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state147_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state147_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state147_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state147_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state147_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state147_66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state147_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state147_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state147_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state147_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state147_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state147_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state147_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state147_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state147_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state147_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state147_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state147_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state147_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state147_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state147_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state147_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state147_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state147_135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state147_135_2 = reservoir_state[135] <<< 2;
wire signed [31:0] shifted_state147_135_3 = reservoir_state[135] <<< 3;
wire signed [31:0] shifted_state147_135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state147_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state147_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state147_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state147_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state147_147_1 = reservoir_state[147] <<< 1;
wire signed [31:0] shifted_state147_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state147_147_5 = reservoir_state[147] <<< 5;
wire signed [31:0] shifted_state147_147_6 = reservoir_state[147] <<< 6;
wire signed [31:0] shifted_state147_147_7 = reservoir_state[147] <<< 7;
wire signed [31:0] shifted_state147_160_1 = reservoir_state[160] <<< 1;
wire signed [31:0] shifted_state147_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state147_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state147_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state147_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state147_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state147_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state147_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state147_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state147_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state147_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state147_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state147_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state147_183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state147_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state147_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state147_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state147_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state147_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state147_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state148_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state148_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state148_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state148_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state148_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state148_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state148_23_0 = reservoir_state[23] <<< 0;
wire signed [31:0] shifted_state148_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state148_23_4 = reservoir_state[23] <<< 4;
wire signed [31:0] shifted_state148_23_5 = reservoir_state[23] <<< 5;
wire signed [31:0] shifted_state148_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state148_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state148_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state148_36_1 = reservoir_state[36] <<< 1;
wire signed [31:0] shifted_state148_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state148_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state148_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state148_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state148_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state148_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state148_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state148_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state148_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state148_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state148_51_6 = reservoir_state[51] <<< 6;
wire signed [31:0] shifted_state148_51_7 = reservoir_state[51] <<< 7;
wire signed [31:0] shifted_state148_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state148_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state148_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state148_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state148_54_4 = reservoir_state[54] <<< 4;
wire signed [31:0] shifted_state148_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state148_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state148_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state148_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state148_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state148_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state148_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state148_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state148_75_3 = reservoir_state[75] <<< 3;
wire signed [31:0] shifted_state148_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state148_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state148_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state148_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state148_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state148_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state148_114_1 = reservoir_state[114] <<< 1;
wire signed [31:0] shifted_state148_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state148_114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state148_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state148_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state148_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state148_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state148_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state148_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state148_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state148_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state148_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state148_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state148_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state148_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state148_169_0 = reservoir_state[169] <<< 0;
wire signed [31:0] shifted_state148_169_2 = reservoir_state[169] <<< 2;
wire signed [31:0] shifted_state148_169_3 = reservoir_state[169] <<< 3;
wire signed [31:0] shifted_state148_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state148_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state148_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state148_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state148_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state148_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state148_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state148_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state148_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state148_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state148_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state148_199_2 = reservoir_state[199] <<< 2;
wire signed [31:0] shifted_state148_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state148_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state148_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state148_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state149_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state149_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state149_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state149_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state149_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state149_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state149_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state149_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state149_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state149_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state149_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state149_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state149_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state149_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state149_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state149_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state149_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state149_103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state149_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state149_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state149_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state149_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state149_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state149_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state149_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state149_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state149_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state149_149_2 = reservoir_state[149] <<< 2;
wire signed [31:0] shifted_state149_149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state149_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state149_149_6 = reservoir_state[149] <<< 6;
wire signed [31:0] shifted_state149_149_7 = reservoir_state[149] <<< 7;
wire signed [31:0] shifted_state149_159_0 = reservoir_state[159] <<< 0;
wire signed [31:0] shifted_state149_159_4 = reservoir_state[159] <<< 4;
wire signed [31:0] shifted_state149_159_5 = reservoir_state[159] <<< 5;
wire signed [31:0] shifted_state149_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state149_160_1 = reservoir_state[160] <<< 1;
wire signed [31:0] shifted_state149_160_2 = reservoir_state[160] <<< 2;
wire signed [31:0] shifted_state149_160_4 = reservoir_state[160] <<< 4;
wire signed [31:0] shifted_state149_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state149_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state149_166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state149_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state149_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state149_167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state149_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state149_167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state149_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state149_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state149_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state149_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state149_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state149_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state149_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state149_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state149_174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state149_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state150_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state150_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state150_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state150_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state150_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state150_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state150_12_2 = reservoir_state[12] <<< 2;
wire signed [31:0] shifted_state150_12_3 = reservoir_state[12] <<< 3;
wire signed [31:0] shifted_state150_12_5 = reservoir_state[12] <<< 5;
wire signed [31:0] shifted_state150_12_6 = reservoir_state[12] <<< 6;
wire signed [31:0] shifted_state150_12_7 = reservoir_state[12] <<< 7;
wire signed [31:0] shifted_state150_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state150_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state150_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state150_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state150_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state150_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state150_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state150_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state150_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state150_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state150_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state150_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state150_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state150_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state150_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state150_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state150_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state150_54_4 = reservoir_state[54] <<< 4;
wire signed [31:0] shifted_state150_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state150_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state150_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state150_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state150_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state150_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state150_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state150_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state150_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state150_60_4 = reservoir_state[60] <<< 4;
wire signed [31:0] shifted_state150_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state150_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state150_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state150_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state150_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state150_68_0 = reservoir_state[68] <<< 0;
wire signed [31:0] shifted_state150_68_2 = reservoir_state[68] <<< 2;
wire signed [31:0] shifted_state150_68_5 = reservoir_state[68] <<< 5;
wire signed [31:0] shifted_state150_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state150_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state150_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state150_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state150_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state150_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state150_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state150_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state150_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state150_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state150_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state150_129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state150_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state150_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state150_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state150_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state150_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state150_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state150_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state150_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state150_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state150_136_3 = reservoir_state[136] <<< 3;
wire signed [31:0] shifted_state150_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state150_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state150_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state150_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state150_148_4 = reservoir_state[148] <<< 4;
wire signed [31:0] shifted_state150_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state150_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state150_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state150_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state150_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state150_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state150_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state150_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state150_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state150_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state150_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state150_170_1 = reservoir_state[170] <<< 1;
wire signed [31:0] shifted_state150_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state150_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state150_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state150_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state150_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state150_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state150_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state150_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state150_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state150_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state150_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state151_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state151_6_3 = reservoir_state[6] <<< 3;
wire signed [31:0] shifted_state151_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state151_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state151_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state151_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state151_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state151_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state151_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state151_18_3 = reservoir_state[18] <<< 3;
wire signed [31:0] shifted_state151_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state151_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state151_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state151_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state151_62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state151_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state151_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state151_62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state151_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state151_62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state151_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state151_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state151_92_4 = reservoir_state[92] <<< 4;
wire signed [31:0] shifted_state151_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state151_92_6 = reservoir_state[92] <<< 6;
wire signed [31:0] shifted_state151_92_7 = reservoir_state[92] <<< 7;
wire signed [31:0] shifted_state151_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state151_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state151_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state151_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state151_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state151_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state151_115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state151_115_6 = reservoir_state[115] <<< 6;
wire signed [31:0] shifted_state151_115_7 = reservoir_state[115] <<< 7;
wire signed [31:0] shifted_state151_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state151_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state151_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state151_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state151_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state151_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state151_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state151_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state151_124_2 = reservoir_state[124] <<< 2;
wire signed [31:0] shifted_state151_124_3 = reservoir_state[124] <<< 3;
wire signed [31:0] shifted_state151_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state151_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state151_124_6 = reservoir_state[124] <<< 6;
wire signed [31:0] shifted_state151_124_7 = reservoir_state[124] <<< 7;
wire signed [31:0] shifted_state151_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state151_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state151_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state151_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state151_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state151_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state151_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state151_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state151_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state151_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state151_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state151_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state151_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state151_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state151_157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state151_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state151_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state151_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state151_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state151_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state151_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state151_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state151_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state151_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state151_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state151_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state152_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state152_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state152_5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state152_5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state152_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state152_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state152_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state152_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state152_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state152_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state152_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state152_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state152_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state152_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state152_35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state152_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state152_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state152_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state152_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state152_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state152_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state152_47_4 = reservoir_state[47] <<< 4;
wire signed [31:0] shifted_state152_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state152_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state152_52_0 = reservoir_state[52] <<< 0;
wire signed [31:0] shifted_state152_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state152_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state152_66_2 = reservoir_state[66] <<< 2;
wire signed [31:0] shifted_state152_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state152_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state152_72_2 = reservoir_state[72] <<< 2;
wire signed [31:0] shifted_state152_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state152_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state152_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state152_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state152_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state152_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state152_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state152_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state152_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state152_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state152_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state152_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state152_90_0 = reservoir_state[90] <<< 0;
wire signed [31:0] shifted_state152_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state152_100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state152_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state152_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state152_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state152_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state152_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state152_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state152_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state152_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state152_102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state152_102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state152_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state152_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state152_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state152_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state152_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state152_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state152_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state152_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state152_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state152_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state152_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state152_139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state152_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state152_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state152_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state152_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state152_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state152_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state153_15_1 = reservoir_state[15] <<< 1;
wire signed [31:0] shifted_state153_15_5 = reservoir_state[15] <<< 5;
wire signed [31:0] shifted_state153_15_6 = reservoir_state[15] <<< 6;
wire signed [31:0] shifted_state153_15_7 = reservoir_state[15] <<< 7;
wire signed [31:0] shifted_state153_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state153_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state153_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state153_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state153_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state153_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state153_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state153_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state153_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state153_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state153_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state153_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state153_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state153_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state153_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state153_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state153_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state153_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state153_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state153_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state153_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state153_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state153_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state153_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state153_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state153_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state153_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state153_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state153_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state153_73_3 = reservoir_state[73] <<< 3;
wire signed [31:0] shifted_state153_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state153_73_5 = reservoir_state[73] <<< 5;
wire signed [31:0] shifted_state153_73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state153_73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state153_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state153_75_4 = reservoir_state[75] <<< 4;
wire signed [31:0] shifted_state153_75_5 = reservoir_state[75] <<< 5;
wire signed [31:0] shifted_state153_75_6 = reservoir_state[75] <<< 6;
wire signed [31:0] shifted_state153_75_7 = reservoir_state[75] <<< 7;
wire signed [31:0] shifted_state153_91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state153_91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state153_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state153_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state153_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state153_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state153_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state153_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state153_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state153_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state153_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state153_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state153_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state153_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state153_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state153_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state153_108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state153_108_4 = reservoir_state[108] <<< 4;
wire signed [31:0] shifted_state153_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state153_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state153_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state153_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state153_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state153_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state153_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state153_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state153_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state153_113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state153_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state153_122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state153_129_0 = reservoir_state[129] <<< 0;
wire signed [31:0] shifted_state153_129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state153_129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state153_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state153_129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state153_129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state153_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state153_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state153_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state153_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state153_140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state153_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state153_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state153_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state153_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state153_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state153_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state153_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state153_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state153_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state153_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state153_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state153_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state153_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state153_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state153_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state153_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state153_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state153_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state153_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state153_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state153_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state153_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state153_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state153_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state153_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state153_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state153_184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state153_184_2 = reservoir_state[184] <<< 2;
wire signed [31:0] shifted_state153_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state153_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state153_184_6 = reservoir_state[184] <<< 6;
wire signed [31:0] shifted_state153_184_7 = reservoir_state[184] <<< 7;
wire signed [31:0] shifted_state154_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state154_8_1 = reservoir_state[8] <<< 1;
wire signed [31:0] shifted_state154_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state154_8_3 = reservoir_state[8] <<< 3;
wire signed [31:0] shifted_state154_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state154_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state154_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state154_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state154_37_2 = reservoir_state[37] <<< 2;
wire signed [31:0] shifted_state154_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state154_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state154_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state154_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state154_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state154_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state154_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state154_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state154_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state154_53_3 = reservoir_state[53] <<< 3;
wire signed [31:0] shifted_state154_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state154_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state154_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state154_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state154_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state154_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state154_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state154_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state154_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state154_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state154_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state154_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state154_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state154_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state154_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state154_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state154_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state154_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state154_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state154_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state154_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state154_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state154_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state154_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state154_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state154_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state154_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state154_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state154_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state154_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state154_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state154_114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state154_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state154_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state154_125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state154_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state154_125_2 = reservoir_state[125] <<< 2;
wire signed [31:0] shifted_state154_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state154_125_5 = reservoir_state[125] <<< 5;
wire signed [31:0] shifted_state154_125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state154_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state154_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state154_157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state154_171_5 = reservoir_state[171] <<< 5;
wire signed [31:0] shifted_state154_171_6 = reservoir_state[171] <<< 6;
wire signed [31:0] shifted_state154_171_7 = reservoir_state[171] <<< 7;
wire signed [31:0] shifted_state154_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state154_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state154_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state154_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state154_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state154_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state154_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state154_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state154_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state154_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state154_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state154_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state154_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state155_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state155_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state155_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state155_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state155_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state155_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state155_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state155_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state155_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state155_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state155_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state155_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state155_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state155_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state155_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state155_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state155_16_3 = reservoir_state[16] <<< 3;
wire signed [31:0] shifted_state155_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state155_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state155_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state155_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state155_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state155_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state155_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state155_60_3 = reservoir_state[60] <<< 3;
wire signed [31:0] shifted_state155_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state155_61_1 = reservoir_state[61] <<< 1;
wire signed [31:0] shifted_state155_61_3 = reservoir_state[61] <<< 3;
wire signed [31:0] shifted_state155_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state155_61_5 = reservoir_state[61] <<< 5;
wire signed [31:0] shifted_state155_61_6 = reservoir_state[61] <<< 6;
wire signed [31:0] shifted_state155_61_7 = reservoir_state[61] <<< 7;
wire signed [31:0] shifted_state155_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state155_72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state155_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state155_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state155_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state155_92_1 = reservoir_state[92] <<< 1;
wire signed [31:0] shifted_state155_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state155_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state155_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state155_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state155_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state155_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state155_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state155_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state155_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state155_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state155_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state155_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state155_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state155_125_5 = reservoir_state[125] <<< 5;
wire signed [31:0] shifted_state155_125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state155_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state155_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state155_131_4 = reservoir_state[131] <<< 4;
wire signed [31:0] shifted_state155_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state155_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state155_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state155_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state155_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state155_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state155_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state155_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state155_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state155_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state155_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state155_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state155_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state155_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state155_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state155_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state155_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state155_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state155_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state155_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state155_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state155_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state155_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state155_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state155_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state155_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state155_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state155_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state155_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state155_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state155_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state155_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state155_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state155_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state155_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state155_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state155_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state155_194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state155_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state155_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state155_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state155_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state156_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state156_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state156_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state156_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state156_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state156_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state156_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state156_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state156_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state156_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state156_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state156_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state156_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state156_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state156_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state156_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state156_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state156_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state156_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state156_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state156_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state156_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state156_38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state156_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state156_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state156_38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state156_40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state156_40_2 = reservoir_state[40] <<< 2;
wire signed [31:0] shifted_state156_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state156_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state156_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state156_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state156_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state156_43_1 = reservoir_state[43] <<< 1;
wire signed [31:0] shifted_state156_43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state156_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state156_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state156_44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state156_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state156_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state156_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state156_44_5 = reservoir_state[44] <<< 5;
wire signed [31:0] shifted_state156_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state156_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state156_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state156_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state156_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state156_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state156_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state156_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state156_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state156_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state156_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state156_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state156_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state156_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state156_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state156_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state156_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state156_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state156_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state156_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state156_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state156_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state156_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state156_168_3 = reservoir_state[168] <<< 3;
wire signed [31:0] shifted_state156_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state156_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state156_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state156_177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state156_177_3 = reservoir_state[177] <<< 3;
wire signed [31:0] shifted_state156_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state156_177_5 = reservoir_state[177] <<< 5;
wire signed [31:0] shifted_state156_177_6 = reservoir_state[177] <<< 6;
wire signed [31:0] shifted_state156_177_7 = reservoir_state[177] <<< 7;
wire signed [31:0] shifted_state156_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state156_183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state156_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state156_183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state156_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state156_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state156_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state156_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state156_194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state156_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state156_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state156_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state156_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state156_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state156_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state156_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state156_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state156_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state156_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state156_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state156_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state156_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state157_9_1 = reservoir_state[9] <<< 1;
wire signed [31:0] shifted_state157_9_5 = reservoir_state[9] <<< 5;
wire signed [31:0] shifted_state157_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state157_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state157_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state157_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state157_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state157_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state157_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state157_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state157_30_4 = reservoir_state[30] <<< 4;
wire signed [31:0] shifted_state157_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state157_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state157_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state157_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state157_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state157_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state157_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state157_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state157_50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state157_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state157_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state157_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state157_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state157_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state157_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state157_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state157_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state157_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state157_87_1 = reservoir_state[87] <<< 1;
wire signed [31:0] shifted_state157_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state157_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state157_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state157_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state157_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state157_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state157_103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state157_103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state157_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state157_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state157_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state157_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state157_117_5 = reservoir_state[117] <<< 5;
wire signed [31:0] shifted_state157_117_6 = reservoir_state[117] <<< 6;
wire signed [31:0] shifted_state157_117_7 = reservoir_state[117] <<< 7;
wire signed [31:0] shifted_state157_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state157_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state157_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state157_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state157_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state157_135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state157_135_2 = reservoir_state[135] <<< 2;
wire signed [31:0] shifted_state157_154_0 = reservoir_state[154] <<< 0;
wire signed [31:0] shifted_state157_154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state157_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state157_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state157_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state157_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state157_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state157_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state158_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state158_3_3 = reservoir_state[3] <<< 3;
wire signed [31:0] shifted_state158_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state158_3_5 = reservoir_state[3] <<< 5;
wire signed [31:0] shifted_state158_3_6 = reservoir_state[3] <<< 6;
wire signed [31:0] shifted_state158_3_7 = reservoir_state[3] <<< 7;
wire signed [31:0] shifted_state158_15_2 = reservoir_state[15] <<< 2;
wire signed [31:0] shifted_state158_15_5 = reservoir_state[15] <<< 5;
wire signed [31:0] shifted_state158_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state158_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state158_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state158_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state158_25_6 = reservoir_state[25] <<< 6;
wire signed [31:0] shifted_state158_25_7 = reservoir_state[25] <<< 7;
wire signed [31:0] shifted_state158_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state158_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state158_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state158_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state158_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state158_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state158_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state158_58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state158_58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state158_58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state158_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state158_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state158_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state158_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state158_67_1 = reservoir_state[67] <<< 1;
wire signed [31:0] shifted_state158_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state158_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state158_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state158_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state158_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state158_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state158_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state158_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state158_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state158_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state158_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state158_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state158_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state158_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state158_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state158_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state158_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state158_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state158_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state158_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state158_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state158_114_1 = reservoir_state[114] <<< 1;
wire signed [31:0] shifted_state158_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state158_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state158_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state158_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state158_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state158_160_4 = reservoir_state[160] <<< 4;
wire signed [31:0] shifted_state158_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state158_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state158_171_0 = reservoir_state[171] <<< 0;
wire signed [31:0] shifted_state158_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state158_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state158_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state158_177_4 = reservoir_state[177] <<< 4;
wire signed [31:0] shifted_state158_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state158_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state158_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state158_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state158_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state158_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state158_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state158_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state158_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state158_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state158_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state159_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state159_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state159_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state159_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state159_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state159_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state159_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state159_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state159_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state159_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state159_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state159_21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state159_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state159_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state159_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state159_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state159_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state159_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state159_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state159_51_6 = reservoir_state[51] <<< 6;
wire signed [31:0] shifted_state159_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state159_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state159_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state159_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state159_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state159_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state159_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state159_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state159_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state159_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state159_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state159_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state159_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state159_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state159_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state159_146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state159_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state159_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state159_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state159_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state159_146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state159_154_0 = reservoir_state[154] <<< 0;
wire signed [31:0] shifted_state159_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state159_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state159_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state159_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state159_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state159_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state159_182_2 = reservoir_state[182] <<< 2;
wire signed [31:0] shifted_state159_182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state159_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state159_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state159_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state159_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state160_16_1 = reservoir_state[16] <<< 1;
wire signed [31:0] shifted_state160_16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state160_16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state160_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state160_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state160_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state160_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state160_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state160_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state160_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state160_33_4 = reservoir_state[33] <<< 4;
wire signed [31:0] shifted_state160_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state160_47_3 = reservoir_state[47] <<< 3;
wire signed [31:0] shifted_state160_47_4 = reservoir_state[47] <<< 4;
wire signed [31:0] shifted_state160_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state160_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state160_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state160_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state160_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state160_56_3 = reservoir_state[56] <<< 3;
wire signed [31:0] shifted_state160_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state160_56_5 = reservoir_state[56] <<< 5;
wire signed [31:0] shifted_state160_56_6 = reservoir_state[56] <<< 6;
wire signed [31:0] shifted_state160_56_7 = reservoir_state[56] <<< 7;
wire signed [31:0] shifted_state160_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state160_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state160_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state160_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state160_69_2 = reservoir_state[69] <<< 2;
wire signed [31:0] shifted_state160_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state160_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state160_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state160_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state160_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state160_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state160_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state160_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state160_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state160_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state160_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state160_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state160_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state160_103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state160_103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state160_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state160_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state160_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state160_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state160_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state160_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state160_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state160_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state160_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state160_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state160_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state160_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state160_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state160_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state160_117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state160_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state160_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state160_118_3 = reservoir_state[118] <<< 3;
wire signed [31:0] shifted_state160_119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state160_124_3 = reservoir_state[124] <<< 3;
wire signed [31:0] shifted_state160_157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state160_157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state160_157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state160_157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state160_157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state160_157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state160_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state160_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state160_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state160_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state160_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state160_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state160_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state160_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state160_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state161_27_0 = reservoir_state[27] <<< 0;
wire signed [31:0] shifted_state161_27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state161_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state161_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state161_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state161_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state161_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state161_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state161_48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state161_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state161_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state161_48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state161_65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state161_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state161_65_3 = reservoir_state[65] <<< 3;
wire signed [31:0] shifted_state161_65_4 = reservoir_state[65] <<< 4;
wire signed [31:0] shifted_state161_65_5 = reservoir_state[65] <<< 5;
wire signed [31:0] shifted_state161_65_6 = reservoir_state[65] <<< 6;
wire signed [31:0] shifted_state161_65_7 = reservoir_state[65] <<< 7;
wire signed [31:0] shifted_state161_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state161_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state161_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state161_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state161_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state161_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state161_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state161_85_7 = reservoir_state[85] <<< 7;
wire signed [31:0] shifted_state161_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state161_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state161_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state161_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state161_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state161_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state161_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state161_111_4 = reservoir_state[111] <<< 4;
wire signed [31:0] shifted_state161_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state161_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state161_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state161_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state161_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state161_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state161_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state161_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state161_113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state161_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state161_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state161_124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state161_124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state161_124_7 = reservoir_state[124] <<< 7;
wire signed [31:0] shifted_state161_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state161_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state161_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state161_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state161_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state161_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state161_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state161_152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state161_152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state161_152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state161_161_0 = reservoir_state[161] <<< 0;
wire signed [31:0] shifted_state161_161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state161_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state161_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state161_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state161_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state161_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state162_9_3 = reservoir_state[9] <<< 3;
wire signed [31:0] shifted_state162_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state162_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state162_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state162_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state162_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state162_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state162_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state162_21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state162_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state162_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state162_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state162_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state162_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state162_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state162_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state162_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state162_25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state162_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state162_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state162_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state162_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state162_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state162_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state162_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state162_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state162_40_2 = reservoir_state[40] <<< 2;
wire signed [31:0] shifted_state162_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state162_40_4 = reservoir_state[40] <<< 4;
wire signed [31:0] shifted_state162_40_5 = reservoir_state[40] <<< 5;
wire signed [31:0] shifted_state162_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state162_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state162_55_2 = reservoir_state[55] <<< 2;
wire signed [31:0] shifted_state162_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state162_55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state162_55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state162_55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state162_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state162_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state162_58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state162_59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state162_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state162_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state162_92_4 = reservoir_state[92] <<< 4;
wire signed [31:0] shifted_state162_92_5 = reservoir_state[92] <<< 5;
wire signed [31:0] shifted_state162_96_1 = reservoir_state[96] <<< 1;
wire signed [31:0] shifted_state162_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state162_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state162_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state162_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state162_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state162_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state162_102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state162_102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state162_102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state162_102_7 = reservoir_state[102] <<< 7;
wire signed [31:0] shifted_state162_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state162_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state162_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state162_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state162_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state162_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state162_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state162_143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state162_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state162_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state162_149_0 = reservoir_state[149] <<< 0;
wire signed [31:0] shifted_state162_149_1 = reservoir_state[149] <<< 1;
wire signed [31:0] shifted_state162_149_4 = reservoir_state[149] <<< 4;
wire signed [31:0] shifted_state162_149_5 = reservoir_state[149] <<< 5;
wire signed [31:0] shifted_state162_149_6 = reservoir_state[149] <<< 6;
wire signed [31:0] shifted_state162_149_7 = reservoir_state[149] <<< 7;
wire signed [31:0] shifted_state162_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state162_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state163_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state163_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state163_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state163_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state163_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state163_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state163_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state163_52_0 = reservoir_state[52] <<< 0;
wire signed [31:0] shifted_state163_52_1 = reservoir_state[52] <<< 1;
wire signed [31:0] shifted_state163_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state163_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state163_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state163_71_0 = reservoir_state[71] <<< 0;
wire signed [31:0] shifted_state163_71_3 = reservoir_state[71] <<< 3;
wire signed [31:0] shifted_state163_71_4 = reservoir_state[71] <<< 4;
wire signed [31:0] shifted_state163_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state163_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state163_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state163_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state163_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state163_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state163_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state163_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state163_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state163_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state163_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state163_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state163_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state163_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state163_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state163_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state163_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state163_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state163_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state163_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state163_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state163_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state163_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state163_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state163_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state163_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state163_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state163_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state163_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state163_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state163_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state163_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state163_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state163_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state163_182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state163_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state163_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state163_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state163_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state163_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state163_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state163_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state163_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state163_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state163_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state163_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state163_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state163_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state163_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state163_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state163_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state163_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state163_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state163_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state163_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state163_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state163_196_4 = reservoir_state[196] <<< 4;
wire signed [31:0] shifted_state163_196_5 = reservoir_state[196] <<< 5;
wire signed [31:0] shifted_state163_196_6 = reservoir_state[196] <<< 6;
wire signed [31:0] shifted_state163_196_7 = reservoir_state[196] <<< 7;
wire signed [31:0] shifted_state163_197_0 = reservoir_state[197] <<< 0;
wire signed [31:0] shifted_state163_197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state163_197_4 = reservoir_state[197] <<< 4;
wire signed [31:0] shifted_state164_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state164_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state164_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state164_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state164_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state164_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state164_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state164_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state164_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state164_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state164_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state164_13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state164_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state164_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state164_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state164_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state164_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state164_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state164_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state164_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state164_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state164_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state164_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state164_29_0 = reservoir_state[29] <<< 0;
wire signed [31:0] shifted_state164_29_4 = reservoir_state[29] <<< 4;
wire signed [31:0] shifted_state164_29_5 = reservoir_state[29] <<< 5;
wire signed [31:0] shifted_state164_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state164_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state164_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state164_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state164_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state164_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state164_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state164_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state164_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state164_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state164_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state164_47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state164_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state164_47_2 = reservoir_state[47] <<< 2;
wire signed [31:0] shifted_state164_47_4 = reservoir_state[47] <<< 4;
wire signed [31:0] shifted_state164_47_5 = reservoir_state[47] <<< 5;
wire signed [31:0] shifted_state164_47_6 = reservoir_state[47] <<< 6;
wire signed [31:0] shifted_state164_47_7 = reservoir_state[47] <<< 7;
wire signed [31:0] shifted_state164_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state164_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state164_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state164_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state164_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state164_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state164_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state164_69_2 = reservoir_state[69] <<< 2;
wire signed [31:0] shifted_state164_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state164_69_5 = reservoir_state[69] <<< 5;
wire signed [31:0] shifted_state164_69_6 = reservoir_state[69] <<< 6;
wire signed [31:0] shifted_state164_69_7 = reservoir_state[69] <<< 7;
wire signed [31:0] shifted_state164_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state164_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state164_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state164_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state164_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state164_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state164_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state164_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state164_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state164_85_2 = reservoir_state[85] <<< 2;
wire signed [31:0] shifted_state164_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state164_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state164_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state164_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state164_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state164_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state164_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state164_94_0 = reservoir_state[94] <<< 0;
wire signed [31:0] shifted_state164_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state164_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state164_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state164_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state164_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state164_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state164_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state164_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state164_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state164_122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state164_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state164_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state164_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state164_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state164_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state164_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state164_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state164_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state164_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state164_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state164_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state164_140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state164_154_0 = reservoir_state[154] <<< 0;
wire signed [31:0] shifted_state164_154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state164_154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state164_154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state164_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state164_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state164_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state164_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state164_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state164_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state164_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state164_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state164_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state164_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state164_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state164_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state164_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state164_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state164_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state164_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state164_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state164_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state164_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state165_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state165_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state165_13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state165_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state165_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state165_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state165_27_0 = reservoir_state[27] <<< 0;
wire signed [31:0] shifted_state165_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state165_27_4 = reservoir_state[27] <<< 4;
wire signed [31:0] shifted_state165_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state165_75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state165_75_1 = reservoir_state[75] <<< 1;
wire signed [31:0] shifted_state165_75_2 = reservoir_state[75] <<< 2;
wire signed [31:0] shifted_state165_75_3 = reservoir_state[75] <<< 3;
wire signed [31:0] shifted_state165_75_4 = reservoir_state[75] <<< 4;
wire signed [31:0] shifted_state165_75_6 = reservoir_state[75] <<< 6;
wire signed [31:0] shifted_state165_75_7 = reservoir_state[75] <<< 7;
wire signed [31:0] shifted_state165_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state165_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state165_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state165_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state165_101_3 = reservoir_state[101] <<< 3;
wire signed [31:0] shifted_state165_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state165_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state165_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state165_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state165_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state165_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state165_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state165_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state165_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state165_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state165_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state165_126_3 = reservoir_state[126] <<< 3;
wire signed [31:0] shifted_state165_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state165_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state165_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state165_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state165_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state165_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state165_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state165_138_0 = reservoir_state[138] <<< 0;
wire signed [31:0] shifted_state165_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state165_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state165_153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state165_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state165_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state165_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state165_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state165_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state165_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state165_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state165_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state165_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state165_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state165_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state165_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state165_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state165_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state165_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state165_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state165_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state166_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state166_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state166_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state166_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state166_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state166_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state166_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state166_3_2 = reservoir_state[3] <<< 2;
wire signed [31:0] shifted_state166_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state166_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state166_16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state166_16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state166_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state166_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state166_17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state166_17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state166_17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state166_26_0 = reservoir_state[26] <<< 0;
wire signed [31:0] shifted_state166_26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state166_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state166_26_5 = reservoir_state[26] <<< 5;
wire signed [31:0] shifted_state166_26_6 = reservoir_state[26] <<< 6;
wire signed [31:0] shifted_state166_26_7 = reservoir_state[26] <<< 7;
wire signed [31:0] shifted_state166_29_3 = reservoir_state[29] <<< 3;
wire signed [31:0] shifted_state166_29_5 = reservoir_state[29] <<< 5;
wire signed [31:0] shifted_state166_29_6 = reservoir_state[29] <<< 6;
wire signed [31:0] shifted_state166_29_7 = reservoir_state[29] <<< 7;
wire signed [31:0] shifted_state166_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state166_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state166_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state166_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state166_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state166_32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state166_32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state166_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state166_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state166_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state166_38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state166_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state166_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state166_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state166_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state166_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state166_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state166_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state166_46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state166_46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state166_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state166_50_5 = reservoir_state[50] <<< 5;
wire signed [31:0] shifted_state166_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state166_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state166_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state166_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state166_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state166_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state166_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state166_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state166_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state166_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state166_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state166_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state166_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state166_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state166_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state166_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state166_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state166_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state166_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state166_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state166_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state166_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state166_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state166_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state166_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state166_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state166_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state166_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state166_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state166_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state166_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state166_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state166_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state166_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state166_158_3 = reservoir_state[158] <<< 3;
wire signed [31:0] shifted_state166_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state166_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state166_158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state166_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state166_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state166_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state166_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state166_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state166_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state166_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state166_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state166_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state166_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state166_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state166_191_0 = reservoir_state[191] <<< 0;
wire signed [31:0] shifted_state166_191_2 = reservoir_state[191] <<< 2;
wire signed [31:0] shifted_state166_191_4 = reservoir_state[191] <<< 4;
wire signed [31:0] shifted_state166_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state166_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state166_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state167_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state167_6_3 = reservoir_state[6] <<< 3;
wire signed [31:0] shifted_state167_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state167_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state167_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state167_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state167_12_0 = reservoir_state[12] <<< 0;
wire signed [31:0] shifted_state167_12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state167_12_2 = reservoir_state[12] <<< 2;
wire signed [31:0] shifted_state167_12_5 = reservoir_state[12] <<< 5;
wire signed [31:0] shifted_state167_12_6 = reservoir_state[12] <<< 6;
wire signed [31:0] shifted_state167_12_7 = reservoir_state[12] <<< 7;
wire signed [31:0] shifted_state167_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state167_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state167_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state167_25_0 = reservoir_state[25] <<< 0;
wire signed [31:0] shifted_state167_25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state167_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state167_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state167_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state167_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state167_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state167_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state167_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state167_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state167_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state167_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state167_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state167_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state167_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state167_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state167_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state167_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state167_57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state167_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state167_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state167_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state167_61_2 = reservoir_state[61] <<< 2;
wire signed [31:0] shifted_state167_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state167_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state167_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state167_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state167_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state167_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state167_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state167_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state167_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state167_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state167_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state167_96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state167_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state167_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state167_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state167_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state167_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state167_103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state167_103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state167_103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state167_106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state167_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state167_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state167_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state167_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state167_107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state167_107_2 = reservoir_state[107] <<< 2;
wire signed [31:0] shifted_state167_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state167_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state167_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state167_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state167_111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state167_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state167_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state167_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state167_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state167_121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state167_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state167_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state167_153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state167_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state167_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state167_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state167_153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state167_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state167_162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state167_162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state167_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state167_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state167_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state167_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state167_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state167_174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state167_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state167_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state167_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state167_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state167_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state167_180_4 = reservoir_state[180] <<< 4;
wire signed [31:0] shifted_state167_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state167_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state167_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state167_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state167_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state167_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state167_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state167_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state167_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state167_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state167_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state167_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state167_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state167_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state168_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state168_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state168_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state168_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state168_19_1 = reservoir_state[19] <<< 1;
wire signed [31:0] shifted_state168_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state168_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state168_20_0 = reservoir_state[20] <<< 0;
wire signed [31:0] shifted_state168_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state168_20_3 = reservoir_state[20] <<< 3;
wire signed [31:0] shifted_state168_20_4 = reservoir_state[20] <<< 4;
wire signed [31:0] shifted_state168_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state168_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state168_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state168_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state168_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state168_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state168_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state168_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state168_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state168_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state168_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state168_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state168_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state168_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state168_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state168_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state168_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state168_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state168_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state168_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state168_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state168_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state168_56_0 = reservoir_state[56] <<< 0;
wire signed [31:0] shifted_state168_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state168_56_4 = reservoir_state[56] <<< 4;
wire signed [31:0] shifted_state168_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state168_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state168_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state168_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state168_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state168_68_1 = reservoir_state[68] <<< 1;
wire signed [31:0] shifted_state168_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state168_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state168_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state168_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state168_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state168_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state168_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state168_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state168_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state168_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state168_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state168_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state168_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state168_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state168_177_0 = reservoir_state[177] <<< 0;
wire signed [31:0] shifted_state168_177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state168_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state168_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state168_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state168_180_5 = reservoir_state[180] <<< 5;
wire signed [31:0] shifted_state168_180_6 = reservoir_state[180] <<< 6;
wire signed [31:0] shifted_state168_180_7 = reservoir_state[180] <<< 7;
wire signed [31:0] shifted_state169_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state169_5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state169_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state169_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state169_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state169_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state169_34_3 = reservoir_state[34] <<< 3;
wire signed [31:0] shifted_state169_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state169_34_6 = reservoir_state[34] <<< 6;
wire signed [31:0] shifted_state169_34_7 = reservoir_state[34] <<< 7;
wire signed [31:0] shifted_state169_50_0 = reservoir_state[50] <<< 0;
wire signed [31:0] shifted_state169_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state169_53_1 = reservoir_state[53] <<< 1;
wire signed [31:0] shifted_state169_53_4 = reservoir_state[53] <<< 4;
wire signed [31:0] shifted_state169_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state169_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state169_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state169_54_5 = reservoir_state[54] <<< 5;
wire signed [31:0] shifted_state169_54_6 = reservoir_state[54] <<< 6;
wire signed [31:0] shifted_state169_54_7 = reservoir_state[54] <<< 7;
wire signed [31:0] shifted_state169_58_1 = reservoir_state[58] <<< 1;
wire signed [31:0] shifted_state169_58_2 = reservoir_state[58] <<< 2;
wire signed [31:0] shifted_state169_77_0 = reservoir_state[77] <<< 0;
wire signed [31:0] shifted_state169_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state169_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state169_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state169_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state169_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state169_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state169_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state169_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state169_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state169_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state169_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state169_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state169_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state169_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state169_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state169_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state169_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state169_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state169_111_2 = reservoir_state[111] <<< 2;
wire signed [31:0] shifted_state169_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state169_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state169_126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state169_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state169_126_3 = reservoir_state[126] <<< 3;
wire signed [31:0] shifted_state169_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state169_129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state169_129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state169_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state169_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state169_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state169_148_4 = reservoir_state[148] <<< 4;
wire signed [31:0] shifted_state169_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state169_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state169_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state169_174_0 = reservoir_state[174] <<< 0;
wire signed [31:0] shifted_state169_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state170_12_0 = reservoir_state[12] <<< 0;
wire signed [31:0] shifted_state170_12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state170_12_5 = reservoir_state[12] <<< 5;
wire signed [31:0] shifted_state170_12_6 = reservoir_state[12] <<< 6;
wire signed [31:0] shifted_state170_12_7 = reservoir_state[12] <<< 7;
wire signed [31:0] shifted_state170_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state170_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state170_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state170_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state170_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state170_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state170_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state170_34_1 = reservoir_state[34] <<< 1;
wire signed [31:0] shifted_state170_34_2 = reservoir_state[34] <<< 2;
wire signed [31:0] shifted_state170_34_5 = reservoir_state[34] <<< 5;
wire signed [31:0] shifted_state170_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state170_66_2 = reservoir_state[66] <<< 2;
wire signed [31:0] shifted_state170_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state170_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state170_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state170_70_2 = reservoir_state[70] <<< 2;
wire signed [31:0] shifted_state170_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state170_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state170_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state170_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state170_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state170_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state170_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state170_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state170_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state170_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state170_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state170_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state170_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state170_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state170_98_5 = reservoir_state[98] <<< 5;
wire signed [31:0] shifted_state170_98_6 = reservoir_state[98] <<< 6;
wire signed [31:0] shifted_state170_98_7 = reservoir_state[98] <<< 7;
wire signed [31:0] shifted_state170_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state170_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state170_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state170_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state170_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state170_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state170_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state170_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state170_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state170_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state170_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state170_124_0 = reservoir_state[124] <<< 0;
wire signed [31:0] shifted_state170_124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state170_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state170_133_2 = reservoir_state[133] <<< 2;
wire signed [31:0] shifted_state170_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state170_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state170_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state170_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state170_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state170_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state170_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state170_162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state170_162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state170_162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state170_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state170_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state170_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state170_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state170_173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state170_173_3 = reservoir_state[173] <<< 3;
wire signed [31:0] shifted_state170_173_4 = reservoir_state[173] <<< 4;
wire signed [31:0] shifted_state170_173_5 = reservoir_state[173] <<< 5;
wire signed [31:0] shifted_state170_173_6 = reservoir_state[173] <<< 6;
wire signed [31:0] shifted_state170_173_7 = reservoir_state[173] <<< 7;
wire signed [31:0] shifted_state171_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state171_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state171_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state171_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state171_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state171_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state171_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state171_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state171_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state171_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state171_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state171_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state171_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state171_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state171_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state171_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state171_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state171_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state171_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state171_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state171_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state171_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state171_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state171_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state171_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state171_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state171_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state171_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state171_83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state171_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state171_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state171_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state171_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state171_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state171_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state171_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state171_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state171_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state171_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state171_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state171_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state171_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state171_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state171_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state171_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state171_139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state171_139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state171_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state171_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state171_139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state171_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state171_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state171_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state171_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state171_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state171_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state171_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state171_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state171_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state171_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state172_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state172_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state172_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state172_5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state172_5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state172_5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state172_5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state172_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state172_8_4 = reservoir_state[8] <<< 4;
wire signed [31:0] shifted_state172_8_5 = reservoir_state[8] <<< 5;
wire signed [31:0] shifted_state172_8_6 = reservoir_state[8] <<< 6;
wire signed [31:0] shifted_state172_8_7 = reservoir_state[8] <<< 7;
wire signed [31:0] shifted_state172_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state172_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state172_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state172_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state172_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state172_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state172_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state172_32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state172_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state172_32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state172_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state172_54_0 = reservoir_state[54] <<< 0;
wire signed [31:0] shifted_state172_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state172_54_2 = reservoir_state[54] <<< 2;
wire signed [31:0] shifted_state172_54_3 = reservoir_state[54] <<< 3;
wire signed [31:0] shifted_state172_54_4 = reservoir_state[54] <<< 4;
wire signed [31:0] shifted_state172_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state172_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state172_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state172_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state172_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state172_72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state172_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state172_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state172_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state172_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state172_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state172_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state172_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state172_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state172_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state172_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state172_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state172_112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state172_119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state172_119_3 = reservoir_state[119] <<< 3;
wire signed [31:0] shifted_state172_119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state172_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state172_128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state172_128_3 = reservoir_state[128] <<< 3;
wire signed [31:0] shifted_state172_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state172_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state172_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state172_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state172_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state172_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state172_134_5 = reservoir_state[134] <<< 5;
wire signed [31:0] shifted_state172_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state172_134_7 = reservoir_state[134] <<< 7;
wire signed [31:0] shifted_state172_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state172_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state172_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state172_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state172_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state172_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state172_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state172_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state172_175_2 = reservoir_state[175] <<< 2;
wire signed [31:0] shifted_state172_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state172_175_4 = reservoir_state[175] <<< 4;
wire signed [31:0] shifted_state172_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state172_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state172_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state172_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state172_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state172_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state172_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state173_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state173_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state173_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state173_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state173_24_3 = reservoir_state[24] <<< 3;
wire signed [31:0] shifted_state173_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state173_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state173_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state173_28_1 = reservoir_state[28] <<< 1;
wire signed [31:0] shifted_state173_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state173_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state173_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state173_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state173_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state173_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state173_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state173_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state173_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state173_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state173_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state173_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state173_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state173_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state173_55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state173_55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state173_55_2 = reservoir_state[55] <<< 2;
wire signed [31:0] shifted_state173_55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state173_55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state173_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state173_58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state173_58_2 = reservoir_state[58] <<< 2;
wire signed [31:0] shifted_state173_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state173_58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state173_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state173_78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state173_78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state173_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state173_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state173_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state173_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state173_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state173_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state173_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state173_110_3 = reservoir_state[110] <<< 3;
wire signed [31:0] shifted_state173_110_4 = reservoir_state[110] <<< 4;
wire signed [31:0] shifted_state173_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state173_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state173_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state173_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state173_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state173_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state173_114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state173_114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state173_153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state173_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state173_153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state173_153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state174_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state174_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state174_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state174_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state174_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state174_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state174_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state174_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state174_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state174_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state174_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state174_57_3 = reservoir_state[57] <<< 3;
wire signed [31:0] shifted_state174_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state174_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state174_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state174_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state174_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state174_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state174_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state174_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state174_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state174_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state174_64_4 = reservoir_state[64] <<< 4;
wire signed [31:0] shifted_state174_79_0 = reservoir_state[79] <<< 0;
wire signed [31:0] shifted_state174_79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state174_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state174_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state174_88_3 = reservoir_state[88] <<< 3;
wire signed [31:0] shifted_state174_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state174_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state174_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state174_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state174_113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state174_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state174_115_3 = reservoir_state[115] <<< 3;
wire signed [31:0] shifted_state174_115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state174_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state174_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state174_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state174_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state174_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state174_145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state174_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state174_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state174_148_4 = reservoir_state[148] <<< 4;
wire signed [31:0] shifted_state174_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state174_151_4 = reservoir_state[151] <<< 4;
wire signed [31:0] shifted_state174_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state174_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state174_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state174_154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state174_154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state174_154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state174_154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state174_154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state174_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state174_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state174_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state174_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state174_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state174_166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state174_166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state174_166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state174_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state174_170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state174_170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state174_170_3 = reservoir_state[170] <<< 3;
wire signed [31:0] shifted_state174_170_4 = reservoir_state[170] <<< 4;
wire signed [31:0] shifted_state174_170_5 = reservoir_state[170] <<< 5;
wire signed [31:0] shifted_state174_170_6 = reservoir_state[170] <<< 6;
wire signed [31:0] shifted_state174_170_7 = reservoir_state[170] <<< 7;
wire signed [31:0] shifted_state174_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state174_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state174_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state174_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state174_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state174_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state174_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state174_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state174_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state174_198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state174_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state174_198_2 = reservoir_state[198] <<< 2;
wire signed [31:0] shifted_state174_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state175_12_3 = reservoir_state[12] <<< 3;
wire signed [31:0] shifted_state175_12_4 = reservoir_state[12] <<< 4;
wire signed [31:0] shifted_state175_12_6 = reservoir_state[12] <<< 6;
wire signed [31:0] shifted_state175_12_7 = reservoir_state[12] <<< 7;
wire signed [31:0] shifted_state175_17_0 = reservoir_state[17] <<< 0;
wire signed [31:0] shifted_state175_17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state175_17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state175_17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state175_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state175_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state175_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state175_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state175_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state175_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state175_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state175_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state175_31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state175_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state175_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state175_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state175_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state175_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state175_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state175_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state175_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state175_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state175_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state175_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state175_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state175_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state175_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state175_68_2 = reservoir_state[68] <<< 2;
wire signed [31:0] shifted_state175_68_3 = reservoir_state[68] <<< 3;
wire signed [31:0] shifted_state175_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state175_69_2 = reservoir_state[69] <<< 2;
wire signed [31:0] shifted_state175_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state175_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state175_69_5 = reservoir_state[69] <<< 5;
wire signed [31:0] shifted_state175_69_6 = reservoir_state[69] <<< 6;
wire signed [31:0] shifted_state175_69_7 = reservoir_state[69] <<< 7;
wire signed [31:0] shifted_state175_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state175_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state175_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state175_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state175_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state175_113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state175_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state175_113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state175_113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state175_120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state175_120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state175_120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state175_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state175_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state175_123_2 = reservoir_state[123] <<< 2;
wire signed [31:0] shifted_state175_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state175_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state175_139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state175_139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state175_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state175_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state175_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state175_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state175_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state175_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state175_176_3 = reservoir_state[176] <<< 3;
wire signed [31:0] shifted_state175_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state175_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state175_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state175_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state175_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state175_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state175_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state175_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state175_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state175_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state176_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state176_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state176_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state176_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state176_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state176_38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state176_38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state176_70_0 = reservoir_state[70] <<< 0;
wire signed [31:0] shifted_state176_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state176_70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state176_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state176_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state176_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state176_79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state176_79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state176_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state176_94_2 = reservoir_state[94] <<< 2;
wire signed [31:0] shifted_state176_94_3 = reservoir_state[94] <<< 3;
wire signed [31:0] shifted_state176_94_4 = reservoir_state[94] <<< 4;
wire signed [31:0] shifted_state176_94_5 = reservoir_state[94] <<< 5;
wire signed [31:0] shifted_state176_94_6 = reservoir_state[94] <<< 6;
wire signed [31:0] shifted_state176_94_7 = reservoir_state[94] <<< 7;
wire signed [31:0] shifted_state176_110_0 = reservoir_state[110] <<< 0;
wire signed [31:0] shifted_state176_110_1 = reservoir_state[110] <<< 1;
wire signed [31:0] shifted_state176_110_3 = reservoir_state[110] <<< 3;
wire signed [31:0] shifted_state176_115_0 = reservoir_state[115] <<< 0;
wire signed [31:0] shifted_state176_115_2 = reservoir_state[115] <<< 2;
wire signed [31:0] shifted_state176_115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state176_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state176_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state176_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state176_130_5 = reservoir_state[130] <<< 5;
wire signed [31:0] shifted_state176_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state176_140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state176_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state176_140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state176_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state176_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state176_144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state176_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state176_144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state176_144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state176_146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state176_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state176_146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state176_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state176_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state176_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state176_148_5 = reservoir_state[148] <<< 5;
wire signed [31:0] shifted_state176_148_6 = reservoir_state[148] <<< 6;
wire signed [31:0] shifted_state176_148_7 = reservoir_state[148] <<< 7;
wire signed [31:0] shifted_state176_173_0 = reservoir_state[173] <<< 0;
wire signed [31:0] shifted_state177_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state177_13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state177_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state177_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state177_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state177_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state177_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state177_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state177_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state177_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state177_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state177_27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state177_27_3 = reservoir_state[27] <<< 3;
wire signed [31:0] shifted_state177_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state177_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state177_30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state177_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state177_30_4 = reservoir_state[30] <<< 4;
wire signed [31:0] shifted_state177_43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state177_43_1 = reservoir_state[43] <<< 1;
wire signed [31:0] shifted_state177_43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state177_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state177_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state177_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state177_67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state177_67_2 = reservoir_state[67] <<< 2;
wire signed [31:0] shifted_state177_67_3 = reservoir_state[67] <<< 3;
wire signed [31:0] shifted_state177_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state177_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state177_76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state177_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state177_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state177_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state177_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state177_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state177_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state177_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state177_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state177_85_3 = reservoir_state[85] <<< 3;
wire signed [31:0] shifted_state177_85_4 = reservoir_state[85] <<< 4;
wire signed [31:0] shifted_state177_85_5 = reservoir_state[85] <<< 5;
wire signed [31:0] shifted_state177_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state177_85_7 = reservoir_state[85] <<< 7;
wire signed [31:0] shifted_state177_138_1 = reservoir_state[138] <<< 1;
wire signed [31:0] shifted_state177_138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state177_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state177_148_0 = reservoir_state[148] <<< 0;
wire signed [31:0] shifted_state177_148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state177_148_2 = reservoir_state[148] <<< 2;
wire signed [31:0] shifted_state177_148_3 = reservoir_state[148] <<< 3;
wire signed [31:0] shifted_state177_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state177_165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state177_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state177_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state177_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state177_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state177_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state177_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state177_172_7 = reservoir_state[172] <<< 7;
wire signed [31:0] shifted_state177_174_1 = reservoir_state[174] <<< 1;
wire signed [31:0] shifted_state177_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state177_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state177_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state177_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state177_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state177_195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state177_198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state177_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state177_198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state177_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state177_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state178_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state178_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state178_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state178_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state178_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state178_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state178_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state178_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state178_21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state178_21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state178_60_0 = reservoir_state[60] <<< 0;
wire signed [31:0] shifted_state178_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state178_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state178_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state178_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state178_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state178_61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state178_61_4 = reservoir_state[61] <<< 4;
wire signed [31:0] shifted_state178_82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state178_82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state178_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state178_82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state178_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state178_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state178_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state178_87_1 = reservoir_state[87] <<< 1;
wire signed [31:0] shifted_state178_87_2 = reservoir_state[87] <<< 2;
wire signed [31:0] shifted_state178_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state178_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state178_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state178_92_1 = reservoir_state[92] <<< 1;
wire signed [31:0] shifted_state178_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state178_92_3 = reservoir_state[92] <<< 3;
wire signed [31:0] shifted_state178_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state178_93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state178_93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state178_93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state178_110_0 = reservoir_state[110] <<< 0;
wire signed [31:0] shifted_state178_110_2 = reservoir_state[110] <<< 2;
wire signed [31:0] shifted_state178_110_3 = reservoir_state[110] <<< 3;
wire signed [31:0] shifted_state178_133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state178_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state178_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state178_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state178_133_6 = reservoir_state[133] <<< 6;
wire signed [31:0] shifted_state178_133_7 = reservoir_state[133] <<< 7;
wire signed [31:0] shifted_state178_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state178_138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state178_138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state178_138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state178_138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state178_144_0 = reservoir_state[144] <<< 0;
wire signed [31:0] shifted_state178_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state178_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state178_144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state178_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state178_164_1 = reservoir_state[164] <<< 1;
wire signed [31:0] shifted_state178_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state178_164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state178_164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state178_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state179_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state179_5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state179_5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state179_5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state179_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state179_6_3 = reservoir_state[6] <<< 3;
wire signed [31:0] shifted_state179_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state179_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state179_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state179_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state179_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state179_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state179_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state179_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state179_20_5 = reservoir_state[20] <<< 5;
wire signed [31:0] shifted_state179_20_6 = reservoir_state[20] <<< 6;
wire signed [31:0] shifted_state179_20_7 = reservoir_state[20] <<< 7;
wire signed [31:0] shifted_state179_22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state179_22_3 = reservoir_state[22] <<< 3;
wire signed [31:0] shifted_state179_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state179_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state179_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state179_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state179_39_0 = reservoir_state[39] <<< 0;
wire signed [31:0] shifted_state179_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state179_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state179_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state179_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state179_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state179_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state179_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state179_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state179_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state179_57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state179_57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state179_57_4 = reservoir_state[57] <<< 4;
wire signed [31:0] shifted_state179_57_5 = reservoir_state[57] <<< 5;
wire signed [31:0] shifted_state179_57_6 = reservoir_state[57] <<< 6;
wire signed [31:0] shifted_state179_57_7 = reservoir_state[57] <<< 7;
wire signed [31:0] shifted_state179_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state179_62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state179_62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state179_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state179_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state179_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state179_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state179_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state179_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state179_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state179_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state179_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state179_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state179_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state179_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state179_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state179_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state179_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state179_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state179_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state179_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state179_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state179_109_0 = reservoir_state[109] <<< 0;
wire signed [31:0] shifted_state179_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state179_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state179_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state179_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state179_111_3 = reservoir_state[111] <<< 3;
wire signed [31:0] shifted_state179_111_5 = reservoir_state[111] <<< 5;
wire signed [31:0] shifted_state179_111_6 = reservoir_state[111] <<< 6;
wire signed [31:0] shifted_state179_111_7 = reservoir_state[111] <<< 7;
wire signed [31:0] shifted_state179_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state179_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state179_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state179_122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state179_122_1 = reservoir_state[122] <<< 1;
wire signed [31:0] shifted_state179_122_3 = reservoir_state[122] <<< 3;
wire signed [31:0] shifted_state179_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state179_122_6 = reservoir_state[122] <<< 6;
wire signed [31:0] shifted_state179_122_7 = reservoir_state[122] <<< 7;
wire signed [31:0] shifted_state179_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state179_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state179_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state179_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state179_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state179_146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state179_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state179_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state179_156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state179_171_0 = reservoir_state[171] <<< 0;
wire signed [31:0] shifted_state179_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state179_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state179_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state179_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state179_193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state179_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state179_193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state179_193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state180_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state180_0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state180_0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state180_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state180_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state180_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state180_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state180_3_0 = reservoir_state[3] <<< 0;
wire signed [31:0] shifted_state180_3_1 = reservoir_state[3] <<< 1;
wire signed [31:0] shifted_state180_3_4 = reservoir_state[3] <<< 4;
wire signed [31:0] shifted_state180_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state180_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state180_18_3 = reservoir_state[18] <<< 3;
wire signed [31:0] shifted_state180_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state180_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state180_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state180_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state180_32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state180_32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state180_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state180_33_0 = reservoir_state[33] <<< 0;
wire signed [31:0] shifted_state180_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state180_33_4 = reservoir_state[33] <<< 4;
wire signed [31:0] shifted_state180_38_0 = reservoir_state[38] <<< 0;
wire signed [31:0] shifted_state180_38_2 = reservoir_state[38] <<< 2;
wire signed [31:0] shifted_state180_38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state180_39_0 = reservoir_state[39] <<< 0;
wire signed [31:0] shifted_state180_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state180_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state180_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state180_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state180_39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state180_39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state180_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state180_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state180_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state180_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state180_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state180_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state180_42_5 = reservoir_state[42] <<< 5;
wire signed [31:0] shifted_state180_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state180_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state180_49_1 = reservoir_state[49] <<< 1;
wire signed [31:0] shifted_state180_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state180_49_3 = reservoir_state[49] <<< 3;
wire signed [31:0] shifted_state180_49_4 = reservoir_state[49] <<< 4;
wire signed [31:0] shifted_state180_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state180_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state180_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state180_66_0 = reservoir_state[66] <<< 0;
wire signed [31:0] shifted_state180_66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state180_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state180_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state180_66_5 = reservoir_state[66] <<< 5;
wire signed [31:0] shifted_state180_66_6 = reservoir_state[66] <<< 6;
wire signed [31:0] shifted_state180_66_7 = reservoir_state[66] <<< 7;
wire signed [31:0] shifted_state180_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state180_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state180_73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state180_73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state180_76_0 = reservoir_state[76] <<< 0;
wire signed [31:0] shifted_state180_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state180_76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state180_76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state180_76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state180_76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state180_77_1 = reservoir_state[77] <<< 1;
wire signed [31:0] shifted_state180_77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state180_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state180_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state180_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state180_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state180_86_1 = reservoir_state[86] <<< 1;
wire signed [31:0] shifted_state180_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state180_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state180_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state180_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state180_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state180_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state180_99_1 = reservoir_state[99] <<< 1;
wire signed [31:0] shifted_state180_99_2 = reservoir_state[99] <<< 2;
wire signed [31:0] shifted_state180_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state180_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state180_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state180_112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state180_112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state180_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state180_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state180_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state180_113_2 = reservoir_state[113] <<< 2;
wire signed [31:0] shifted_state180_113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state180_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state180_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state180_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state180_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state180_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state180_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state180_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state180_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state180_143_2 = reservoir_state[143] <<< 2;
wire signed [31:0] shifted_state180_143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state180_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state180_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state180_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state180_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state180_145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state180_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state180_147_3 = reservoir_state[147] <<< 3;
wire signed [31:0] shifted_state180_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state180_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state180_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state180_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state180_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state180_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state180_164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state180_164_2 = reservoir_state[164] <<< 2;
wire signed [31:0] shifted_state180_164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state180_164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state180_164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state180_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state180_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state180_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state180_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state180_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state180_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state180_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state180_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state180_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state180_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state180_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state180_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state180_193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state180_193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state181_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state181_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state181_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state181_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state181_23_1 = reservoir_state[23] <<< 1;
wire signed [31:0] shifted_state181_23_2 = reservoir_state[23] <<< 2;
wire signed [31:0] shifted_state181_23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state181_23_5 = reservoir_state[23] <<< 5;
wire signed [31:0] shifted_state181_23_6 = reservoir_state[23] <<< 6;
wire signed [31:0] shifted_state181_23_7 = reservoir_state[23] <<< 7;
wire signed [31:0] shifted_state181_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state181_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state181_28_5 = reservoir_state[28] <<< 5;
wire signed [31:0] shifted_state181_28_6 = reservoir_state[28] <<< 6;
wire signed [31:0] shifted_state181_28_7 = reservoir_state[28] <<< 7;
wire signed [31:0] shifted_state181_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state181_35_3 = reservoir_state[35] <<< 3;
wire signed [31:0] shifted_state181_35_4 = reservoir_state[35] <<< 4;
wire signed [31:0] shifted_state181_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state181_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state181_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state181_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state181_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state181_37_5 = reservoir_state[37] <<< 5;
wire signed [31:0] shifted_state181_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state181_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state181_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state181_46_1 = reservoir_state[46] <<< 1;
wire signed [31:0] shifted_state181_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state181_46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state181_53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state181_53_5 = reservoir_state[53] <<< 5;
wire signed [31:0] shifted_state181_53_6 = reservoir_state[53] <<< 6;
wire signed [31:0] shifted_state181_53_7 = reservoir_state[53] <<< 7;
wire signed [31:0] shifted_state181_67_2 = reservoir_state[67] <<< 2;
wire signed [31:0] shifted_state181_67_5 = reservoir_state[67] <<< 5;
wire signed [31:0] shifted_state181_67_6 = reservoir_state[67] <<< 6;
wire signed [31:0] shifted_state181_67_7 = reservoir_state[67] <<< 7;
wire signed [31:0] shifted_state181_73_1 = reservoir_state[73] <<< 1;
wire signed [31:0] shifted_state181_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state181_74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state181_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state181_74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state181_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state181_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state181_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state181_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state181_80_3 = reservoir_state[80] <<< 3;
wire signed [31:0] shifted_state181_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state181_80_6 = reservoir_state[80] <<< 6;
wire signed [31:0] shifted_state181_80_7 = reservoir_state[80] <<< 7;
wire signed [31:0] shifted_state181_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state181_85_1 = reservoir_state[85] <<< 1;
wire signed [31:0] shifted_state181_85_3 = reservoir_state[85] <<< 3;
wire signed [31:0] shifted_state181_92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state181_92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state181_92_4 = reservoir_state[92] <<< 4;
wire signed [31:0] shifted_state181_92_6 = reservoir_state[92] <<< 6;
wire signed [31:0] shifted_state181_92_7 = reservoir_state[92] <<< 7;
wire signed [31:0] shifted_state181_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state181_104_3 = reservoir_state[104] <<< 3;
wire signed [31:0] shifted_state181_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state181_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state181_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state181_137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state181_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state181_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state181_144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state181_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state181_144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state181_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state181_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state181_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state181_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state181_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state181_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state181_151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state181_151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state181_151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state181_151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state181_151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state181_151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state181_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state181_168_2 = reservoir_state[168] <<< 2;
wire signed [31:0] shifted_state181_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state181_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state181_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state181_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state181_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state181_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state181_190_0 = reservoir_state[190] <<< 0;
wire signed [31:0] shifted_state181_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state181_190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state181_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state181_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state181_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state181_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state182_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state182_27_0 = reservoir_state[27] <<< 0;
wire signed [31:0] shifted_state182_27_6 = reservoir_state[27] <<< 6;
wire signed [31:0] shifted_state182_27_7 = reservoir_state[27] <<< 7;
wire signed [31:0] shifted_state182_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state182_36_4 = reservoir_state[36] <<< 4;
wire signed [31:0] shifted_state182_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state182_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state182_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state182_48_0 = reservoir_state[48] <<< 0;
wire signed [31:0] shifted_state182_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state182_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state182_48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state182_52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state182_52_4 = reservoir_state[52] <<< 4;
wire signed [31:0] shifted_state182_52_5 = reservoir_state[52] <<< 5;
wire signed [31:0] shifted_state182_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state182_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state182_64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state182_64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state182_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state182_65_4 = reservoir_state[65] <<< 4;
wire signed [31:0] shifted_state182_65_5 = reservoir_state[65] <<< 5;
wire signed [31:0] shifted_state182_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state182_93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state182_99_0 = reservoir_state[99] <<< 0;
wire signed [31:0] shifted_state182_99_3 = reservoir_state[99] <<< 3;
wire signed [31:0] shifted_state182_99_4 = reservoir_state[99] <<< 4;
wire signed [31:0] shifted_state182_99_5 = reservoir_state[99] <<< 5;
wire signed [31:0] shifted_state182_99_6 = reservoir_state[99] <<< 6;
wire signed [31:0] shifted_state182_99_7 = reservoir_state[99] <<< 7;
wire signed [31:0] shifted_state182_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state182_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state182_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state182_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state182_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state182_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state182_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state182_175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state182_175_3 = reservoir_state[175] <<< 3;
wire signed [31:0] shifted_state182_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state182_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state182_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state182_178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state182_178_3 = reservoir_state[178] <<< 3;
wire signed [31:0] shifted_state182_178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state182_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state182_185_2 = reservoir_state[185] <<< 2;
wire signed [31:0] shifted_state182_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state182_185_5 = reservoir_state[185] <<< 5;
wire signed [31:0] shifted_state182_185_6 = reservoir_state[185] <<< 6;
wire signed [31:0] shifted_state182_185_7 = reservoir_state[185] <<< 7;
wire signed [31:0] shifted_state182_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state182_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state182_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state182_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state182_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state182_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state182_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state182_197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state182_197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state182_197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state182_197_7 = reservoir_state[197] <<< 7;
wire signed [31:0] shifted_state183_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state183_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state183_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state183_25_2 = reservoir_state[25] <<< 2;
wire signed [31:0] shifted_state183_25_3 = reservoir_state[25] <<< 3;
wire signed [31:0] shifted_state183_25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state183_37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state183_37_3 = reservoir_state[37] <<< 3;
wire signed [31:0] shifted_state183_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state183_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state183_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state183_44_3 = reservoir_state[44] <<< 3;
wire signed [31:0] shifted_state183_52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state183_52_4 = reservoir_state[52] <<< 4;
wire signed [31:0] shifted_state183_52_5 = reservoir_state[52] <<< 5;
wire signed [31:0] shifted_state183_52_6 = reservoir_state[52] <<< 6;
wire signed [31:0] shifted_state183_52_7 = reservoir_state[52] <<< 7;
wire signed [31:0] shifted_state183_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state183_64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state183_64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state183_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state183_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state183_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state183_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state183_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state183_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state183_97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state183_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state183_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state183_110_1 = reservoir_state[110] <<< 1;
wire signed [31:0] shifted_state183_110_3 = reservoir_state[110] <<< 3;
wire signed [31:0] shifted_state183_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state183_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state183_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state183_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state183_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state183_131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state183_131_1 = reservoir_state[131] <<< 1;
wire signed [31:0] shifted_state183_131_2 = reservoir_state[131] <<< 2;
wire signed [31:0] shifted_state183_131_3 = reservoir_state[131] <<< 3;
wire signed [31:0] shifted_state183_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state183_140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state183_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state183_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state183_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state183_144_1 = reservoir_state[144] <<< 1;
wire signed [31:0] shifted_state183_144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state183_144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state183_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state183_161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state183_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state183_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state183_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state183_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state183_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state183_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state183_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state183_165_4 = reservoir_state[165] <<< 4;
wire signed [31:0] shifted_state183_165_5 = reservoir_state[165] <<< 5;
wire signed [31:0] shifted_state183_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state183_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state183_167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state183_167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state183_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state183_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state184_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state184_2_3 = reservoir_state[2] <<< 3;
wire signed [31:0] shifted_state184_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state184_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state184_28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state184_28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state184_28_3 = reservoir_state[28] <<< 3;
wire signed [31:0] shifted_state184_28_4 = reservoir_state[28] <<< 4;
wire signed [31:0] shifted_state184_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state184_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state184_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state184_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state184_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state184_34_4 = reservoir_state[34] <<< 4;
wire signed [31:0] shifted_state184_35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state184_35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state184_35_5 = reservoir_state[35] <<< 5;
wire signed [31:0] shifted_state184_35_6 = reservoir_state[35] <<< 6;
wire signed [31:0] shifted_state184_35_7 = reservoir_state[35] <<< 7;
wire signed [31:0] shifted_state184_37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state184_37_4 = reservoir_state[37] <<< 4;
wire signed [31:0] shifted_state184_37_6 = reservoir_state[37] <<< 6;
wire signed [31:0] shifted_state184_37_7 = reservoir_state[37] <<< 7;
wire signed [31:0] shifted_state184_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state184_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state184_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state184_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state184_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state184_42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state184_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state184_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state184_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state184_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state184_46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state184_46_2 = reservoir_state[46] <<< 2;
wire signed [31:0] shifted_state184_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state184_50_3 = reservoir_state[50] <<< 3;
wire signed [31:0] shifted_state184_52_1 = reservoir_state[52] <<< 1;
wire signed [31:0] shifted_state184_52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state184_52_4 = reservoir_state[52] <<< 4;
wire signed [31:0] shifted_state184_52_5 = reservoir_state[52] <<< 5;
wire signed [31:0] shifted_state184_52_6 = reservoir_state[52] <<< 6;
wire signed [31:0] shifted_state184_52_7 = reservoir_state[52] <<< 7;
wire signed [31:0] shifted_state184_70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state184_70_2 = reservoir_state[70] <<< 2;
wire signed [31:0] shifted_state184_70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state184_70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state184_70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state184_71_2 = reservoir_state[71] <<< 2;
wire signed [31:0] shifted_state184_71_5 = reservoir_state[71] <<< 5;
wire signed [31:0] shifted_state184_71_6 = reservoir_state[71] <<< 6;
wire signed [31:0] shifted_state184_71_7 = reservoir_state[71] <<< 7;
wire signed [31:0] shifted_state184_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state184_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state184_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state184_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state184_101_0 = reservoir_state[101] <<< 0;
wire signed [31:0] shifted_state184_101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state184_101_2 = reservoir_state[101] <<< 2;
wire signed [31:0] shifted_state184_101_3 = reservoir_state[101] <<< 3;
wire signed [31:0] shifted_state184_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state184_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state184_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state184_114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state184_114_1 = reservoir_state[114] <<< 1;
wire signed [31:0] shifted_state184_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state184_114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state184_117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state184_117_1 = reservoir_state[117] <<< 1;
wire signed [31:0] shifted_state184_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state184_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state184_117_6 = reservoir_state[117] <<< 6;
wire signed [31:0] shifted_state184_117_7 = reservoir_state[117] <<< 7;
wire signed [31:0] shifted_state184_134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state184_134_3 = reservoir_state[134] <<< 3;
wire signed [31:0] shifted_state184_134_6 = reservoir_state[134] <<< 6;
wire signed [31:0] shifted_state184_134_7 = reservoir_state[134] <<< 7;
wire signed [31:0] shifted_state184_140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state184_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state184_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state184_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state184_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state184_165_6 = reservoir_state[165] <<< 6;
wire signed [31:0] shifted_state184_165_7 = reservoir_state[165] <<< 7;
wire signed [31:0] shifted_state184_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state184_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state184_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state184_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state184_192_1 = reservoir_state[192] <<< 1;
wire signed [31:0] shifted_state184_192_3 = reservoir_state[192] <<< 3;
wire signed [31:0] shifted_state184_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state184_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state184_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state184_193_1 = reservoir_state[193] <<< 1;
wire signed [31:0] shifted_state184_193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state184_193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state185_2_0 = reservoir_state[2] <<< 0;
wire signed [31:0] shifted_state185_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state185_2_5 = reservoir_state[2] <<< 5;
wire signed [31:0] shifted_state185_2_6 = reservoir_state[2] <<< 6;
wire signed [31:0] shifted_state185_2_7 = reservoir_state[2] <<< 7;
wire signed [31:0] shifted_state185_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state185_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state185_6_3 = reservoir_state[6] <<< 3;
wire signed [31:0] shifted_state185_6_4 = reservoir_state[6] <<< 4;
wire signed [31:0] shifted_state185_6_6 = reservoir_state[6] <<< 6;
wire signed [31:0] shifted_state185_6_7 = reservoir_state[6] <<< 7;
wire signed [31:0] shifted_state185_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state185_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state185_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state185_15_4 = reservoir_state[15] <<< 4;
wire signed [31:0] shifted_state185_15_6 = reservoir_state[15] <<< 6;
wire signed [31:0] shifted_state185_15_7 = reservoir_state[15] <<< 7;
wire signed [31:0] shifted_state185_46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state185_46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state185_47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state185_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state185_49_3 = reservoir_state[49] <<< 3;
wire signed [31:0] shifted_state185_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state185_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state185_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state185_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state185_50_4 = reservoir_state[50] <<< 4;
wire signed [31:0] shifted_state185_50_6 = reservoir_state[50] <<< 6;
wire signed [31:0] shifted_state185_50_7 = reservoir_state[50] <<< 7;
wire signed [31:0] shifted_state185_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state185_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state185_69_4 = reservoir_state[69] <<< 4;
wire signed [31:0] shifted_state185_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state185_87_1 = reservoir_state[87] <<< 1;
wire signed [31:0] shifted_state185_87_2 = reservoir_state[87] <<< 2;
wire signed [31:0] shifted_state185_87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state185_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state185_87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state185_87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state185_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state185_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state185_93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state185_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state185_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state185_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state185_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state185_115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state185_115_4 = reservoir_state[115] <<< 4;
wire signed [31:0] shifted_state185_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state185_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state185_133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state185_133_3 = reservoir_state[133] <<< 3;
wire signed [31:0] shifted_state185_133_4 = reservoir_state[133] <<< 4;
wire signed [31:0] shifted_state185_160_1 = reservoir_state[160] <<< 1;
wire signed [31:0] shifted_state185_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state185_169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state185_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state185_169_5 = reservoir_state[169] <<< 5;
wire signed [31:0] shifted_state185_169_6 = reservoir_state[169] <<< 6;
wire signed [31:0] shifted_state185_169_7 = reservoir_state[169] <<< 7;
wire signed [31:0] shifted_state185_185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state185_185_3 = reservoir_state[185] <<< 3;
wire signed [31:0] shifted_state185_185_4 = reservoir_state[185] <<< 4;
wire signed [31:0] shifted_state186_8_0 = reservoir_state[8] <<< 0;
wire signed [31:0] shifted_state186_8_1 = reservoir_state[8] <<< 1;
wire signed [31:0] shifted_state186_8_2 = reservoir_state[8] <<< 2;
wire signed [31:0] shifted_state186_8_3 = reservoir_state[8] <<< 3;
wire signed [31:0] shifted_state186_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state186_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state186_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state186_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state186_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state186_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state186_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state186_14_4 = reservoir_state[14] <<< 4;
wire signed [31:0] shifted_state186_14_6 = reservoir_state[14] <<< 6;
wire signed [31:0] shifted_state186_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state186_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state186_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state186_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state186_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state186_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state186_45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state186_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state186_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state186_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state186_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state186_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state186_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state186_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state186_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state186_73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state186_73_1 = reservoir_state[73] <<< 1;
wire signed [31:0] shifted_state186_73_2 = reservoir_state[73] <<< 2;
wire signed [31:0] shifted_state186_73_3 = reservoir_state[73] <<< 3;
wire signed [31:0] shifted_state186_73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state186_83_0 = reservoir_state[83] <<< 0;
wire signed [31:0] shifted_state186_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state186_83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state186_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state186_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state186_85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state186_85_6 = reservoir_state[85] <<< 6;
wire signed [31:0] shifted_state186_86_3 = reservoir_state[86] <<< 3;
wire signed [31:0] shifted_state186_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state186_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state186_88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state186_88_1 = reservoir_state[88] <<< 1;
wire signed [31:0] shifted_state186_88_2 = reservoir_state[88] <<< 2;
wire signed [31:0] shifted_state186_88_4 = reservoir_state[88] <<< 4;
wire signed [31:0] shifted_state186_110_0 = reservoir_state[110] <<< 0;
wire signed [31:0] shifted_state186_110_2 = reservoir_state[110] <<< 2;
wire signed [31:0] shifted_state186_110_3 = reservoir_state[110] <<< 3;
wire signed [31:0] shifted_state186_110_5 = reservoir_state[110] <<< 5;
wire signed [31:0] shifted_state186_110_6 = reservoir_state[110] <<< 6;
wire signed [31:0] shifted_state186_110_7 = reservoir_state[110] <<< 7;
wire signed [31:0] shifted_state186_125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state186_125_2 = reservoir_state[125] <<< 2;
wire signed [31:0] shifted_state186_125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state186_125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state186_125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state186_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state186_133_5 = reservoir_state[133] <<< 5;
wire signed [31:0] shifted_state186_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state186_147_1 = reservoir_state[147] <<< 1;
wire signed [31:0] shifted_state186_147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state186_147_3 = reservoir_state[147] <<< 3;
wire signed [31:0] shifted_state186_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state186_153_1 = reservoir_state[153] <<< 1;
wire signed [31:0] shifted_state186_153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state186_153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state186_156_0 = reservoir_state[156] <<< 0;
wire signed [31:0] shifted_state186_156_1 = reservoir_state[156] <<< 1;
wire signed [31:0] shifted_state186_156_2 = reservoir_state[156] <<< 2;
wire signed [31:0] shifted_state186_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state186_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state186_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state186_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state187_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state187_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state187_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state187_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state187_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state187_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state187_12_0 = reservoir_state[12] <<< 0;
wire signed [31:0] shifted_state187_12_2 = reservoir_state[12] <<< 2;
wire signed [31:0] shifted_state187_12_3 = reservoir_state[12] <<< 3;
wire signed [31:0] shifted_state187_12_5 = reservoir_state[12] <<< 5;
wire signed [31:0] shifted_state187_20_1 = reservoir_state[20] <<< 1;
wire signed [31:0] shifted_state187_20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state187_40_0 = reservoir_state[40] <<< 0;
wire signed [31:0] shifted_state187_40_3 = reservoir_state[40] <<< 3;
wire signed [31:0] shifted_state187_40_5 = reservoir_state[40] <<< 5;
wire signed [31:0] shifted_state187_40_6 = reservoir_state[40] <<< 6;
wire signed [31:0] shifted_state187_40_7 = reservoir_state[40] <<< 7;
wire signed [31:0] shifted_state187_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state187_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state187_49_1 = reservoir_state[49] <<< 1;
wire signed [31:0] shifted_state187_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state187_49_6 = reservoir_state[49] <<< 6;
wire signed [31:0] shifted_state187_49_7 = reservoir_state[49] <<< 7;
wire signed [31:0] shifted_state187_58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state187_60_1 = reservoir_state[60] <<< 1;
wire signed [31:0] shifted_state187_60_2 = reservoir_state[60] <<< 2;
wire signed [31:0] shifted_state187_60_4 = reservoir_state[60] <<< 4;
wire signed [31:0] shifted_state187_60_5 = reservoir_state[60] <<< 5;
wire signed [31:0] shifted_state187_60_6 = reservoir_state[60] <<< 6;
wire signed [31:0] shifted_state187_60_7 = reservoir_state[60] <<< 7;
wire signed [31:0] shifted_state187_62_0 = reservoir_state[62] <<< 0;
wire signed [31:0] shifted_state187_62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state187_86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state187_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state187_86_5 = reservoir_state[86] <<< 5;
wire signed [31:0] shifted_state187_86_6 = reservoir_state[86] <<< 6;
wire signed [31:0] shifted_state187_86_7 = reservoir_state[86] <<< 7;
wire signed [31:0] shifted_state187_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state187_97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state187_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state187_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state187_97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state187_97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state187_97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state187_100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state187_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state187_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state187_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state187_100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state187_100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state187_105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state187_105_1 = reservoir_state[105] <<< 1;
wire signed [31:0] shifted_state187_105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state187_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state187_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state187_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state187_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state187_111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state187_137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state187_137_1 = reservoir_state[137] <<< 1;
wire signed [31:0] shifted_state187_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state187_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state187_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state187_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state187_140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state187_140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state187_140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state187_140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state187_140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state187_140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state187_140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state187_147_1 = reservoir_state[147] <<< 1;
wire signed [31:0] shifted_state187_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state187_147_6 = reservoir_state[147] <<< 6;
wire signed [31:0] shifted_state187_147_7 = reservoir_state[147] <<< 7;
wire signed [31:0] shifted_state187_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state187_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state187_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state187_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state187_150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state187_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state187_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state187_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state187_171_3 = reservoir_state[171] <<< 3;
wire signed [31:0] shifted_state187_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state187_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state187_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state187_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state187_183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state187_183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state187_183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state187_183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state187_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state187_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state187_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state187_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state187_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state188_4_1 = reservoir_state[4] <<< 1;
wire signed [31:0] shifted_state188_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state188_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state188_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state188_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state188_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state188_5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state188_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state188_5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state188_5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state188_5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state188_18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state188_18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state188_18_2 = reservoir_state[18] <<< 2;
wire signed [31:0] shifted_state188_18_3 = reservoir_state[18] <<< 3;
wire signed [31:0] shifted_state188_18_4 = reservoir_state[18] <<< 4;
wire signed [31:0] shifted_state188_18_5 = reservoir_state[18] <<< 5;
wire signed [31:0] shifted_state188_18_6 = reservoir_state[18] <<< 6;
wire signed [31:0] shifted_state188_18_7 = reservoir_state[18] <<< 7;
wire signed [31:0] shifted_state188_33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state188_33_2 = reservoir_state[33] <<< 2;
wire signed [31:0] shifted_state188_33_5 = reservoir_state[33] <<< 5;
wire signed [31:0] shifted_state188_33_6 = reservoir_state[33] <<< 6;
wire signed [31:0] shifted_state188_33_7 = reservoir_state[33] <<< 7;
wire signed [31:0] shifted_state188_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state188_42_1 = reservoir_state[42] <<< 1;
wire signed [31:0] shifted_state188_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state188_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state188_42_6 = reservoir_state[42] <<< 6;
wire signed [31:0] shifted_state188_42_7 = reservoir_state[42] <<< 7;
wire signed [31:0] shifted_state188_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state188_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state188_44_6 = reservoir_state[44] <<< 6;
wire signed [31:0] shifted_state188_44_7 = reservoir_state[44] <<< 7;
wire signed [31:0] shifted_state188_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state188_45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state188_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state188_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state188_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state188_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state188_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state188_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state188_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state188_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state188_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state188_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state188_100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state188_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state188_104_5 = reservoir_state[104] <<< 5;
wire signed [31:0] shifted_state188_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state188_104_7 = reservoir_state[104] <<< 7;
wire signed [31:0] shifted_state188_106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state188_106_2 = reservoir_state[106] <<< 2;
wire signed [31:0] shifted_state188_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state188_106_4 = reservoir_state[106] <<< 4;
wire signed [31:0] shifted_state188_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state188_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state188_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state188_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state188_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state188_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state188_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state188_117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state188_117_3 = reservoir_state[117] <<< 3;
wire signed [31:0] shifted_state188_117_4 = reservoir_state[117] <<< 4;
wire signed [31:0] shifted_state188_117_6 = reservoir_state[117] <<< 6;
wire signed [31:0] shifted_state188_117_7 = reservoir_state[117] <<< 7;
wire signed [31:0] shifted_state188_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state188_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state188_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state188_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state188_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state188_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state188_130_4 = reservoir_state[130] <<< 4;
wire signed [31:0] shifted_state188_130_6 = reservoir_state[130] <<< 6;
wire signed [31:0] shifted_state188_130_7 = reservoir_state[130] <<< 7;
wire signed [31:0] shifted_state188_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state188_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state188_142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state188_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state188_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state188_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state188_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state188_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state188_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state188_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state188_155_1 = reservoir_state[155] <<< 1;
wire signed [31:0] shifted_state188_155_2 = reservoir_state[155] <<< 2;
wire signed [31:0] shifted_state188_186_0 = reservoir_state[186] <<< 0;
wire signed [31:0] shifted_state188_186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state188_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state188_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state188_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state188_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state188_192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state188_192_2 = reservoir_state[192] <<< 2;
wire signed [31:0] shifted_state188_192_4 = reservoir_state[192] <<< 4;
wire signed [31:0] shifted_state188_192_5 = reservoir_state[192] <<< 5;
wire signed [31:0] shifted_state188_192_6 = reservoir_state[192] <<< 6;
wire signed [31:0] shifted_state188_192_7 = reservoir_state[192] <<< 7;
wire signed [31:0] shifted_state188_195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state188_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state188_197_2 = reservoir_state[197] <<< 2;
wire signed [31:0] shifted_state188_197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state188_197_4 = reservoir_state[197] <<< 4;
wire signed [31:0] shifted_state188_197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state188_197_7 = reservoir_state[197] <<< 7;
wire signed [31:0] shifted_state189_14_0 = reservoir_state[14] <<< 0;
wire signed [31:0] shifted_state189_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state189_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state189_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state189_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state189_36_0 = reservoir_state[36] <<< 0;
wire signed [31:0] shifted_state189_36_1 = reservoir_state[36] <<< 1;
wire signed [31:0] shifted_state189_36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state189_36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state189_36_4 = reservoir_state[36] <<< 4;
wire signed [31:0] shifted_state189_36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state189_36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state189_36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state189_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state189_39_2 = reservoir_state[39] <<< 2;
wire signed [31:0] shifted_state189_39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state189_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state189_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state189_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state189_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state189_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state189_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state189_48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state189_48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state189_67_1 = reservoir_state[67] <<< 1;
wire signed [31:0] shifted_state189_67_2 = reservoir_state[67] <<< 2;
wire signed [31:0] shifted_state189_67_3 = reservoir_state[67] <<< 3;
wire signed [31:0] shifted_state189_67_4 = reservoir_state[67] <<< 4;
wire signed [31:0] shifted_state189_72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state189_72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state189_72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state189_72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state189_72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state189_78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state189_78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state189_78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state189_78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state189_78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state189_95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state189_95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state189_95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state189_95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state189_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state189_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state189_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state189_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state189_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state189_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state189_130_0 = reservoir_state[130] <<< 0;
wire signed [31:0] shifted_state189_130_1 = reservoir_state[130] <<< 1;
wire signed [31:0] shifted_state189_130_2 = reservoir_state[130] <<< 2;
wire signed [31:0] shifted_state189_130_3 = reservoir_state[130] <<< 3;
wire signed [31:0] shifted_state189_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state189_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state189_141_6 = reservoir_state[141] <<< 6;
wire signed [31:0] shifted_state189_141_7 = reservoir_state[141] <<< 7;
wire signed [31:0] shifted_state189_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state189_150_1 = reservoir_state[150] <<< 1;
wire signed [31:0] shifted_state189_150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state189_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state189_161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state189_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state189_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state189_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state189_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state189_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state189_189_0 = reservoir_state[189] <<< 0;
wire signed [31:0] shifted_state189_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state189_194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state189_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state189_194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state189_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state189_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state189_196_0 = reservoir_state[196] <<< 0;
wire signed [31:0] shifted_state189_196_2 = reservoir_state[196] <<< 2;
wire signed [31:0] shifted_state189_196_3 = reservoir_state[196] <<< 3;
wire signed [31:0] shifted_state189_196_4 = reservoir_state[196] <<< 4;
wire signed [31:0] shifted_state189_196_6 = reservoir_state[196] <<< 6;
wire signed [31:0] shifted_state189_196_7 = reservoir_state[196] <<< 7;
wire signed [31:0] shifted_state190_11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state190_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state190_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state190_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state190_11_5 = reservoir_state[11] <<< 5;
wire signed [31:0] shifted_state190_11_6 = reservoir_state[11] <<< 6;
wire signed [31:0] shifted_state190_11_7 = reservoir_state[11] <<< 7;
wire signed [31:0] shifted_state190_15_3 = reservoir_state[15] <<< 3;
wire signed [31:0] shifted_state190_15_5 = reservoir_state[15] <<< 5;
wire signed [31:0] shifted_state190_15_6 = reservoir_state[15] <<< 6;
wire signed [31:0] shifted_state190_15_7 = reservoir_state[15] <<< 7;
wire signed [31:0] shifted_state190_21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state190_21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state190_21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state190_21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state190_62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state190_65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state190_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state190_65_2 = reservoir_state[65] <<< 2;
wire signed [31:0] shifted_state190_65_5 = reservoir_state[65] <<< 5;
wire signed [31:0] shifted_state190_65_6 = reservoir_state[65] <<< 6;
wire signed [31:0] shifted_state190_65_7 = reservoir_state[65] <<< 7;
wire signed [31:0] shifted_state190_66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state190_66_3 = reservoir_state[66] <<< 3;
wire signed [31:0] shifted_state190_66_4 = reservoir_state[66] <<< 4;
wire signed [31:0] shifted_state190_80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state190_80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state190_80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state190_80_4 = reservoir_state[80] <<< 4;
wire signed [31:0] shifted_state190_80_5 = reservoir_state[80] <<< 5;
wire signed [31:0] shifted_state190_91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state190_91_2 = reservoir_state[91] <<< 2;
wire signed [31:0] shifted_state190_91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state190_91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state190_91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state190_91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state190_97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state190_97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state190_97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state190_107_1 = reservoir_state[107] <<< 1;
wire signed [31:0] shifted_state190_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state190_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state190_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state190_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state190_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state190_109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state190_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state190_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state190_160_0 = reservoir_state[160] <<< 0;
wire signed [31:0] shifted_state190_160_2 = reservoir_state[160] <<< 2;
wire signed [31:0] shifted_state190_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state190_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state190_172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state190_172_2 = reservoir_state[172] <<< 2;
wire signed [31:0] shifted_state190_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state190_172_5 = reservoir_state[172] <<< 5;
wire signed [31:0] shifted_state190_175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state190_175_5 = reservoir_state[175] <<< 5;
wire signed [31:0] shifted_state190_175_6 = reservoir_state[175] <<< 6;
wire signed [31:0] shifted_state190_175_7 = reservoir_state[175] <<< 7;
wire signed [31:0] shifted_state190_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state190_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state190_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state190_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state190_189_6 = reservoir_state[189] <<< 6;
wire signed [31:0] shifted_state190_189_7 = reservoir_state[189] <<< 7;
wire signed [31:0] shifted_state190_194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state190_199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state190_199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state190_199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state190_199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state190_199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state190_199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_state191_1_1 = reservoir_state[1] <<< 1;
wire signed [31:0] shifted_state191_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state191_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state191_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state191_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state191_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state191_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state191_6_3 = reservoir_state[6] <<< 3;
wire signed [31:0] shifted_state191_13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state191_13_1 = reservoir_state[13] <<< 1;
wire signed [31:0] shifted_state191_13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state191_13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state191_13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state191_13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state191_26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state191_26_3 = reservoir_state[26] <<< 3;
wire signed [31:0] shifted_state191_26_4 = reservoir_state[26] <<< 4;
wire signed [31:0] shifted_state191_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state191_30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state191_30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state191_30_4 = reservoir_state[30] <<< 4;
wire signed [31:0] shifted_state191_30_5 = reservoir_state[30] <<< 5;
wire signed [31:0] shifted_state191_30_6 = reservoir_state[30] <<< 6;
wire signed [31:0] shifted_state191_30_7 = reservoir_state[30] <<< 7;
wire signed [31:0] shifted_state191_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state191_43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state191_43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state191_43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state191_45_0 = reservoir_state[45] <<< 0;
wire signed [31:0] shifted_state191_45_1 = reservoir_state[45] <<< 1;
wire signed [31:0] shifted_state191_45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state191_45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state191_45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state191_45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state191_56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state191_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state191_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state191_59_3 = reservoir_state[59] <<< 3;
wire signed [31:0] shifted_state191_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state191_59_5 = reservoir_state[59] <<< 5;
wire signed [31:0] shifted_state191_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state191_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state191_69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state191_69_1 = reservoir_state[69] <<< 1;
wire signed [31:0] shifted_state191_69_3 = reservoir_state[69] <<< 3;
wire signed [31:0] shifted_state191_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state191_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state191_84_2 = reservoir_state[84] <<< 2;
wire signed [31:0] shifted_state191_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state191_98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state191_98_3 = reservoir_state[98] <<< 3;
wire signed [31:0] shifted_state191_98_4 = reservoir_state[98] <<< 4;
wire signed [31:0] shifted_state191_98_5 = reservoir_state[98] <<< 5;
wire signed [31:0] shifted_state191_106_3 = reservoir_state[106] <<< 3;
wire signed [31:0] shifted_state191_106_5 = reservoir_state[106] <<< 5;
wire signed [31:0] shifted_state191_106_6 = reservoir_state[106] <<< 6;
wire signed [31:0] shifted_state191_106_7 = reservoir_state[106] <<< 7;
wire signed [31:0] shifted_state191_132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state191_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state191_132_2 = reservoir_state[132] <<< 2;
wire signed [31:0] shifted_state191_132_4 = reservoir_state[132] <<< 4;
wire signed [31:0] shifted_state191_147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state191_147_4 = reservoir_state[147] <<< 4;
wire signed [31:0] shifted_state191_147_5 = reservoir_state[147] <<< 5;
wire signed [31:0] shifted_state191_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state191_169_4 = reservoir_state[169] <<< 4;
wire signed [31:0] shifted_state191_174_2 = reservoir_state[174] <<< 2;
wire signed [31:0] shifted_state191_174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state191_174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state191_174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state191_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state191_179_2 = reservoir_state[179] <<< 2;
wire signed [31:0] shifted_state191_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state191_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state191_187_0 = reservoir_state[187] <<< 0;
wire signed [31:0] shifted_state191_187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state191_187_2 = reservoir_state[187] <<< 2;
wire signed [31:0] shifted_state191_187_3 = reservoir_state[187] <<< 3;
wire signed [31:0] shifted_state191_187_4 = reservoir_state[187] <<< 4;
wire signed [31:0] shifted_state191_187_5 = reservoir_state[187] <<< 5;
wire signed [31:0] shifted_state191_187_6 = reservoir_state[187] <<< 6;
wire signed [31:0] shifted_state191_187_7 = reservoir_state[187] <<< 7;
wire signed [31:0] shifted_state191_194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state191_194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state191_194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state191_194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state191_194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state191_197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state191_197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state191_197_4 = reservoir_state[197] <<< 4;
wire signed [31:0] shifted_state192_1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state192_1_1 = reservoir_state[1] <<< 1;
wire signed [31:0] shifted_state192_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state192_1_3 = reservoir_state[1] <<< 3;
wire signed [31:0] shifted_state192_1_4 = reservoir_state[1] <<< 4;
wire signed [31:0] shifted_state192_1_5 = reservoir_state[1] <<< 5;
wire signed [31:0] shifted_state192_1_6 = reservoir_state[1] <<< 6;
wire signed [31:0] shifted_state192_1_7 = reservoir_state[1] <<< 7;
wire signed [31:0] shifted_state192_19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state192_19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state192_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state192_19_5 = reservoir_state[19] <<< 5;
wire signed [31:0] shifted_state192_19_6 = reservoir_state[19] <<< 6;
wire signed [31:0] shifted_state192_19_7 = reservoir_state[19] <<< 7;
wire signed [31:0] shifted_state192_22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state192_22_2 = reservoir_state[22] <<< 2;
wire signed [31:0] shifted_state192_22_4 = reservoir_state[22] <<< 4;
wire signed [31:0] shifted_state192_22_5 = reservoir_state[22] <<< 5;
wire signed [31:0] shifted_state192_22_6 = reservoir_state[22] <<< 6;
wire signed [31:0] shifted_state192_22_7 = reservoir_state[22] <<< 7;
wire signed [31:0] shifted_state192_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state192_24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state192_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state192_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state192_24_5 = reservoir_state[24] <<< 5;
wire signed [31:0] shifted_state192_24_6 = reservoir_state[24] <<< 6;
wire signed [31:0] shifted_state192_24_7 = reservoir_state[24] <<< 7;
wire signed [31:0] shifted_state192_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state192_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state192_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state192_44_0 = reservoir_state[44] <<< 0;
wire signed [31:0] shifted_state192_44_2 = reservoir_state[44] <<< 2;
wire signed [31:0] shifted_state192_54_1 = reservoir_state[54] <<< 1;
wire signed [31:0] shifted_state192_54_4 = reservoir_state[54] <<< 4;
wire signed [31:0] shifted_state192_63_0 = reservoir_state[63] <<< 0;
wire signed [31:0] shifted_state192_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state192_63_5 = reservoir_state[63] <<< 5;
wire signed [31:0] shifted_state192_63_6 = reservoir_state[63] <<< 6;
wire signed [31:0] shifted_state192_63_7 = reservoir_state[63] <<< 7;
wire signed [31:0] shifted_state192_77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state192_77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state192_77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state192_77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state192_77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state192_81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state192_81_1 = reservoir_state[81] <<< 1;
wire signed [31:0] shifted_state192_81_3 = reservoir_state[81] <<< 3;
wire signed [31:0] shifted_state192_81_4 = reservoir_state[81] <<< 4;
wire signed [31:0] shifted_state192_81_5 = reservoir_state[81] <<< 5;
wire signed [31:0] shifted_state192_81_6 = reservoir_state[81] <<< 6;
wire signed [31:0] shifted_state192_81_7 = reservoir_state[81] <<< 7;
wire signed [31:0] shifted_state192_93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state192_93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state192_93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state192_93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state192_94_1 = reservoir_state[94] <<< 1;
wire signed [31:0] shifted_state192_94_2 = reservoir_state[94] <<< 2;
wire signed [31:0] shifted_state192_95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state192_95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state192_95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state192_95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state192_96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state192_96_4 = reservoir_state[96] <<< 4;
wire signed [31:0] shifted_state192_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state192_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state192_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state192_103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state192_103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state192_103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state192_103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state192_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state192_112_3 = reservoir_state[112] <<< 3;
wire signed [31:0] shifted_state192_112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state192_112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state192_112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state192_114_2 = reservoir_state[114] <<< 2;
wire signed [31:0] shifted_state192_114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state192_116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state192_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state192_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state192_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state192_118_0 = reservoir_state[118] <<< 0;
wire signed [31:0] shifted_state192_118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state192_118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state192_118_4 = reservoir_state[118] <<< 4;
wire signed [31:0] shifted_state192_118_5 = reservoir_state[118] <<< 5;
wire signed [31:0] shifted_state192_118_6 = reservoir_state[118] <<< 6;
wire signed [31:0] shifted_state192_118_7 = reservoir_state[118] <<< 7;
wire signed [31:0] shifted_state192_123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state192_123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state192_123_3 = reservoir_state[123] <<< 3;
wire signed [31:0] shifted_state192_123_4 = reservoir_state[123] <<< 4;
wire signed [31:0] shifted_state192_123_5 = reservoir_state[123] <<< 5;
wire signed [31:0] shifted_state192_123_6 = reservoir_state[123] <<< 6;
wire signed [31:0] shifted_state192_123_7 = reservoir_state[123] <<< 7;
wire signed [31:0] shifted_state192_136_1 = reservoir_state[136] <<< 1;
wire signed [31:0] shifted_state192_136_2 = reservoir_state[136] <<< 2;
wire signed [31:0] shifted_state192_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state192_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state192_136_6 = reservoir_state[136] <<< 6;
wire signed [31:0] shifted_state192_136_7 = reservoir_state[136] <<< 7;
wire signed [31:0] shifted_state192_161_0 = reservoir_state[161] <<< 0;
wire signed [31:0] shifted_state192_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state192_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state192_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state192_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state192_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state192_166_2 = reservoir_state[166] <<< 2;
wire signed [31:0] shifted_state192_166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state192_166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state192_166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state193_1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state193_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state193_16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state193_16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state193_39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state193_39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state193_39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state193_41_1 = reservoir_state[41] <<< 1;
wire signed [31:0] shifted_state193_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state193_41_3 = reservoir_state[41] <<< 3;
wire signed [31:0] shifted_state193_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state193_41_5 = reservoir_state[41] <<< 5;
wire signed [31:0] shifted_state193_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state193_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state193_50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state193_51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state193_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state193_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state193_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state193_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state193_67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state193_67_1 = reservoir_state[67] <<< 1;
wire signed [31:0] shifted_state193_67_2 = reservoir_state[67] <<< 2;
wire signed [31:0] shifted_state193_67_4 = reservoir_state[67] <<< 4;
wire signed [31:0] shifted_state193_67_6 = reservoir_state[67] <<< 6;
wire signed [31:0] shifted_state193_67_7 = reservoir_state[67] <<< 7;
wire signed [31:0] shifted_state193_84_2 = reservoir_state[84] <<< 2;
wire signed [31:0] shifted_state193_84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state193_86_0 = reservoir_state[86] <<< 0;
wire signed [31:0] shifted_state193_86_4 = reservoir_state[86] <<< 4;
wire signed [31:0] shifted_state193_89_0 = reservoir_state[89] <<< 0;
wire signed [31:0] shifted_state193_89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state193_90_1 = reservoir_state[90] <<< 1;
wire signed [31:0] shifted_state193_90_2 = reservoir_state[90] <<< 2;
wire signed [31:0] shifted_state193_90_6 = reservoir_state[90] <<< 6;
wire signed [31:0] shifted_state193_90_7 = reservoir_state[90] <<< 7;
wire signed [31:0] shifted_state193_100_2 = reservoir_state[100] <<< 2;
wire signed [31:0] shifted_state193_100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state193_100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state193_101_2 = reservoir_state[101] <<< 2;
wire signed [31:0] shifted_state193_101_3 = reservoir_state[101] <<< 3;
wire signed [31:0] shifted_state193_101_4 = reservoir_state[101] <<< 4;
wire signed [31:0] shifted_state193_101_5 = reservoir_state[101] <<< 5;
wire signed [31:0] shifted_state193_101_6 = reservoir_state[101] <<< 6;
wire signed [31:0] shifted_state193_101_7 = reservoir_state[101] <<< 7;
wire signed [31:0] shifted_state193_102_0 = reservoir_state[102] <<< 0;
wire signed [31:0] shifted_state193_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state193_102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state193_102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state193_104_0 = reservoir_state[104] <<< 0;
wire signed [31:0] shifted_state193_104_1 = reservoir_state[104] <<< 1;
wire signed [31:0] shifted_state193_104_2 = reservoir_state[104] <<< 2;
wire signed [31:0] shifted_state193_104_4 = reservoir_state[104] <<< 4;
wire signed [31:0] shifted_state193_104_6 = reservoir_state[104] <<< 6;
wire signed [31:0] shifted_state193_107_3 = reservoir_state[107] <<< 3;
wire signed [31:0] shifted_state193_107_4 = reservoir_state[107] <<< 4;
wire signed [31:0] shifted_state193_107_5 = reservoir_state[107] <<< 5;
wire signed [31:0] shifted_state193_107_6 = reservoir_state[107] <<< 6;
wire signed [31:0] shifted_state193_107_7 = reservoir_state[107] <<< 7;
wire signed [31:0] shifted_state193_108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state193_108_2 = reservoir_state[108] <<< 2;
wire signed [31:0] shifted_state193_108_5 = reservoir_state[108] <<< 5;
wire signed [31:0] shifted_state193_108_6 = reservoir_state[108] <<< 6;
wire signed [31:0] shifted_state193_108_7 = reservoir_state[108] <<< 7;
wire signed [31:0] shifted_state193_113_0 = reservoir_state[113] <<< 0;
wire signed [31:0] shifted_state193_113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state193_113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state193_128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state193_128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state193_128_4 = reservoir_state[128] <<< 4;
wire signed [31:0] shifted_state193_128_5 = reservoir_state[128] <<< 5;
wire signed [31:0] shifted_state193_128_6 = reservoir_state[128] <<< 6;
wire signed [31:0] shifted_state193_128_7 = reservoir_state[128] <<< 7;
wire signed [31:0] shifted_state193_132_1 = reservoir_state[132] <<< 1;
wire signed [31:0] shifted_state193_132_3 = reservoir_state[132] <<< 3;
wire signed [31:0] shifted_state193_132_5 = reservoir_state[132] <<< 5;
wire signed [31:0] shifted_state193_132_6 = reservoir_state[132] <<< 6;
wire signed [31:0] shifted_state193_132_7 = reservoir_state[132] <<< 7;
wire signed [31:0] shifted_state193_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state193_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state193_145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state193_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state193_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state193_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state193_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state193_162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state193_162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state193_162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state193_162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state193_162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state193_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state193_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state193_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state193_168_0 = reservoir_state[168] <<< 0;
wire signed [31:0] shifted_state193_168_1 = reservoir_state[168] <<< 1;
wire signed [31:0] shifted_state193_168_4 = reservoir_state[168] <<< 4;
wire signed [31:0] shifted_state193_168_5 = reservoir_state[168] <<< 5;
wire signed [31:0] shifted_state193_168_6 = reservoir_state[168] <<< 6;
wire signed [31:0] shifted_state193_168_7 = reservoir_state[168] <<< 7;
wire signed [31:0] shifted_state193_181_2 = reservoir_state[181] <<< 2;
wire signed [31:0] shifted_state193_184_3 = reservoir_state[184] <<< 3;
wire signed [31:0] shifted_state193_184_5 = reservoir_state[184] <<< 5;
wire signed [31:0] shifted_state194_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state194_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state194_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state194_30_0 = reservoir_state[30] <<< 0;
wire signed [31:0] shifted_state194_30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state194_30_5 = reservoir_state[30] <<< 5;
wire signed [31:0] shifted_state194_31_0 = reservoir_state[31] <<< 0;
wire signed [31:0] shifted_state194_31_1 = reservoir_state[31] <<< 1;
wire signed [31:0] shifted_state194_31_2 = reservoir_state[31] <<< 2;
wire signed [31:0] shifted_state194_31_4 = reservoir_state[31] <<< 4;
wire signed [31:0] shifted_state194_31_5 = reservoir_state[31] <<< 5;
wire signed [31:0] shifted_state194_31_6 = reservoir_state[31] <<< 6;
wire signed [31:0] shifted_state194_31_7 = reservoir_state[31] <<< 7;
wire signed [31:0] shifted_state194_32_2 = reservoir_state[32] <<< 2;
wire signed [31:0] shifted_state194_32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state194_122_4 = reservoir_state[122] <<< 4;
wire signed [31:0] shifted_state194_122_5 = reservoir_state[122] <<< 5;
wire signed [31:0] shifted_state194_127_0 = reservoir_state[127] <<< 0;
wire signed [31:0] shifted_state194_127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state194_127_2 = reservoir_state[127] <<< 2;
wire signed [31:0] shifted_state194_127_3 = reservoir_state[127] <<< 3;
wire signed [31:0] shifted_state194_127_4 = reservoir_state[127] <<< 4;
wire signed [31:0] shifted_state194_127_5 = reservoir_state[127] <<< 5;
wire signed [31:0] shifted_state194_127_6 = reservoir_state[127] <<< 6;
wire signed [31:0] shifted_state194_127_7 = reservoir_state[127] <<< 7;
wire signed [31:0] shifted_state194_155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state194_155_3 = reservoir_state[155] <<< 3;
wire signed [31:0] shifted_state194_155_4 = reservoir_state[155] <<< 4;
wire signed [31:0] shifted_state194_155_5 = reservoir_state[155] <<< 5;
wire signed [31:0] shifted_state194_155_6 = reservoir_state[155] <<< 6;
wire signed [31:0] shifted_state194_155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state194_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state194_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state194_179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state194_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state194_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state194_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state194_183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state194_183_1 = reservoir_state[183] <<< 1;
wire signed [31:0] shifted_state194_183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state194_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state194_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state194_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state194_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state194_189_5 = reservoir_state[189] <<< 5;
wire signed [31:0] shifted_state194_189_6 = reservoir_state[189] <<< 6;
wire signed [31:0] shifted_state194_189_7 = reservoir_state[189] <<< 7;
wire signed [31:0] shifted_state195_14_0 = reservoir_state[14] <<< 0;
wire signed [31:0] shifted_state195_14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state195_14_2 = reservoir_state[14] <<< 2;
wire signed [31:0] shifted_state195_14_3 = reservoir_state[14] <<< 3;
wire signed [31:0] shifted_state195_14_5 = reservoir_state[14] <<< 5;
wire signed [31:0] shifted_state195_14_7 = reservoir_state[14] <<< 7;
wire signed [31:0] shifted_state195_19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state195_19_4 = reservoir_state[19] <<< 4;
wire signed [31:0] shifted_state195_63_1 = reservoir_state[63] <<< 1;
wire signed [31:0] shifted_state195_63_2 = reservoir_state[63] <<< 2;
wire signed [31:0] shifted_state195_63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state195_63_4 = reservoir_state[63] <<< 4;
wire signed [31:0] shifted_state195_67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state195_67_3 = reservoir_state[67] <<< 3;
wire signed [31:0] shifted_state195_67_6 = reservoir_state[67] <<< 6;
wire signed [31:0] shifted_state195_67_7 = reservoir_state[67] <<< 7;
wire signed [31:0] shifted_state195_74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state195_74_1 = reservoir_state[74] <<< 1;
wire signed [31:0] shifted_state195_96_3 = reservoir_state[96] <<< 3;
wire signed [31:0] shifted_state195_96_5 = reservoir_state[96] <<< 5;
wire signed [31:0] shifted_state195_96_6 = reservoir_state[96] <<< 6;
wire signed [31:0] shifted_state195_96_7 = reservoir_state[96] <<< 7;
wire signed [31:0] shifted_state195_98_0 = reservoir_state[98] <<< 0;
wire signed [31:0] shifted_state195_98_1 = reservoir_state[98] <<< 1;
wire signed [31:0] shifted_state195_109_1 = reservoir_state[109] <<< 1;
wire signed [31:0] shifted_state195_109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state195_109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state195_109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state195_109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state195_109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state195_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state195_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state195_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state195_126_6 = reservoir_state[126] <<< 6;
wire signed [31:0] shifted_state195_126_7 = reservoir_state[126] <<< 7;
wire signed [31:0] shifted_state195_139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state195_139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state195_141_0 = reservoir_state[141] <<< 0;
wire signed [31:0] shifted_state195_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state195_141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state195_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state195_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state195_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state195_145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state195_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state195_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state195_145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state195_145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state195_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state195_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state195_163_3 = reservoir_state[163] <<< 3;
wire signed [31:0] shifted_state195_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state195_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state195_163_6 = reservoir_state[163] <<< 6;
wire signed [31:0] shifted_state195_163_7 = reservoir_state[163] <<< 7;
wire signed [31:0] shifted_state195_171_1 = reservoir_state[171] <<< 1;
wire signed [31:0] shifted_state195_171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state195_171_4 = reservoir_state[171] <<< 4;
wire signed [31:0] shifted_state195_178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state195_178_1 = reservoir_state[178] <<< 1;
wire signed [31:0] shifted_state195_178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state195_178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state195_178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state195_190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state195_190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state195_190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state195_190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state195_190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state195_190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state195_195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state195_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state195_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state195_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state195_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state196_4_0 = reservoir_state[4] <<< 0;
wire signed [31:0] shifted_state196_4_2 = reservoir_state[4] <<< 2;
wire signed [31:0] shifted_state196_4_3 = reservoir_state[4] <<< 3;
wire signed [31:0] shifted_state196_4_4 = reservoir_state[4] <<< 4;
wire signed [31:0] shifted_state196_4_5 = reservoir_state[4] <<< 5;
wire signed [31:0] shifted_state196_4_6 = reservoir_state[4] <<< 6;
wire signed [31:0] shifted_state196_4_7 = reservoir_state[4] <<< 7;
wire signed [31:0] shifted_state196_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state196_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state196_7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state196_7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state196_7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state196_43_1 = reservoir_state[43] <<< 1;
wire signed [31:0] shifted_state196_43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state196_49_0 = reservoir_state[49] <<< 0;
wire signed [31:0] shifted_state196_49_2 = reservoir_state[49] <<< 2;
wire signed [31:0] shifted_state196_49_3 = reservoir_state[49] <<< 3;
wire signed [31:0] shifted_state196_49_5 = reservoir_state[49] <<< 5;
wire signed [31:0] shifted_state196_51_1 = reservoir_state[51] <<< 1;
wire signed [31:0] shifted_state196_51_2 = reservoir_state[51] <<< 2;
wire signed [31:0] shifted_state196_51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state196_51_4 = reservoir_state[51] <<< 4;
wire signed [31:0] shifted_state196_51_5 = reservoir_state[51] <<< 5;
wire signed [31:0] shifted_state196_51_6 = reservoir_state[51] <<< 6;
wire signed [31:0] shifted_state196_51_7 = reservoir_state[51] <<< 7;
wire signed [31:0] shifted_state196_74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state196_74_4 = reservoir_state[74] <<< 4;
wire signed [31:0] shifted_state196_74_5 = reservoir_state[74] <<< 5;
wire signed [31:0] shifted_state196_74_6 = reservoir_state[74] <<< 6;
wire signed [31:0] shifted_state196_74_7 = reservoir_state[74] <<< 7;
wire signed [31:0] shifted_state196_76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state196_76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state196_102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state196_102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state196_112_0 = reservoir_state[112] <<< 0;
wire signed [31:0] shifted_state196_112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state196_112_2 = reservoir_state[112] <<< 2;
wire signed [31:0] shifted_state196_126_0 = reservoir_state[126] <<< 0;
wire signed [31:0] shifted_state196_126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state196_126_4 = reservoir_state[126] <<< 4;
wire signed [31:0] shifted_state196_126_5 = reservoir_state[126] <<< 5;
wire signed [31:0] shifted_state196_142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state196_142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state196_142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state196_142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state196_142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state196_142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state196_165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state196_165_1 = reservoir_state[165] <<< 1;
wire signed [31:0] shifted_state196_165_3 = reservoir_state[165] <<< 3;
wire signed [31:0] shifted_state196_172_0 = reservoir_state[172] <<< 0;
wire signed [31:0] shifted_state196_172_3 = reservoir_state[172] <<< 3;
wire signed [31:0] shifted_state196_172_4 = reservoir_state[172] <<< 4;
wire signed [31:0] shifted_state196_172_6 = reservoir_state[172] <<< 6;
wire signed [31:0] shifted_state196_180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state196_180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state196_180_2 = reservoir_state[180] <<< 2;
wire signed [31:0] shifted_state196_180_3 = reservoir_state[180] <<< 3;
wire signed [31:0] shifted_state196_182_1 = reservoir_state[182] <<< 1;
wire signed [31:0] shifted_state196_182_4 = reservoir_state[182] <<< 4;
wire signed [31:0] shifted_state196_182_5 = reservoir_state[182] <<< 5;
wire signed [31:0] shifted_state196_182_6 = reservoir_state[182] <<< 6;
wire signed [31:0] shifted_state196_182_7 = reservoir_state[182] <<< 7;
wire signed [31:0] shifted_state196_198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state196_198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state196_198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state196_198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state197_0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state197_0_1 = reservoir_state[0] <<< 1;
wire signed [31:0] shifted_state197_0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state197_0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state197_0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state197_0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state197_44_4 = reservoir_state[44] <<< 4;
wire signed [31:0] shifted_state197_87_0 = reservoir_state[87] <<< 0;
wire signed [31:0] shifted_state197_87_2 = reservoir_state[87] <<< 2;
wire signed [31:0] shifted_state197_87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state197_89_1 = reservoir_state[89] <<< 1;
wire signed [31:0] shifted_state197_89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state197_89_4 = reservoir_state[89] <<< 4;
wire signed [31:0] shifted_state197_89_5 = reservoir_state[89] <<< 5;
wire signed [31:0] shifted_state197_89_6 = reservoir_state[89] <<< 6;
wire signed [31:0] shifted_state197_89_7 = reservoir_state[89] <<< 7;
wire signed [31:0] shifted_state197_90_0 = reservoir_state[90] <<< 0;
wire signed [31:0] shifted_state197_90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state197_90_5 = reservoir_state[90] <<< 5;
wire signed [31:0] shifted_state197_121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state197_121_1 = reservoir_state[121] <<< 1;
wire signed [31:0] shifted_state197_121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state197_121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state197_121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state197_121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state197_121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state197_137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state197_137_3 = reservoir_state[137] <<< 3;
wire signed [31:0] shifted_state197_137_4 = reservoir_state[137] <<< 4;
wire signed [31:0] shifted_state197_137_5 = reservoir_state[137] <<< 5;
wire signed [31:0] shifted_state197_137_6 = reservoir_state[137] <<< 6;
wire signed [31:0] shifted_state197_137_7 = reservoir_state[137] <<< 7;
wire signed [31:0] shifted_state197_141_1 = reservoir_state[141] <<< 1;
wire signed [31:0] shifted_state197_141_3 = reservoir_state[141] <<< 3;
wire signed [31:0] shifted_state197_141_4 = reservoir_state[141] <<< 4;
wire signed [31:0] shifted_state197_141_5 = reservoir_state[141] <<< 5;
wire signed [31:0] shifted_state197_143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state197_143_3 = reservoir_state[143] <<< 3;
wire signed [31:0] shifted_state197_143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state197_143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state197_143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state197_143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state197_150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state197_150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state197_150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state197_150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state197_150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state197_152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state197_156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state197_156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state197_156_6 = reservoir_state[156] <<< 6;
wire signed [31:0] shifted_state197_156_7 = reservoir_state[156] <<< 7;
wire signed [31:0] shifted_state197_159_0 = reservoir_state[159] <<< 0;
wire signed [31:0] shifted_state197_159_2 = reservoir_state[159] <<< 2;
wire signed [31:0] shifted_state197_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state197_159_4 = reservoir_state[159] <<< 4;
wire signed [31:0] shifted_state197_159_6 = reservoir_state[159] <<< 6;
wire signed [31:0] shifted_state197_159_7 = reservoir_state[159] <<< 7;
wire signed [31:0] shifted_state197_163_0 = reservoir_state[163] <<< 0;
wire signed [31:0] shifted_state197_163_1 = reservoir_state[163] <<< 1;
wire signed [31:0] shifted_state197_163_2 = reservoir_state[163] <<< 2;
wire signed [31:0] shifted_state197_163_4 = reservoir_state[163] <<< 4;
wire signed [31:0] shifted_state197_163_5 = reservoir_state[163] <<< 5;
wire signed [31:0] shifted_state197_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state197_176_2 = reservoir_state[176] <<< 2;
wire signed [31:0] shifted_state197_176_3 = reservoir_state[176] <<< 3;
wire signed [31:0] shifted_state197_195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state197_195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state197_195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state197_195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state197_195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state198_5_0 = reservoir_state[5] <<< 0;
wire signed [31:0] shifted_state198_5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state198_5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state198_5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state198_5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state198_5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state198_7_0 = reservoir_state[7] <<< 0;
wire signed [31:0] shifted_state198_7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state198_7_2 = reservoir_state[7] <<< 2;
wire signed [31:0] shifted_state198_7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state198_7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state198_9_4 = reservoir_state[9] <<< 4;
wire signed [31:0] shifted_state198_10_0 = reservoir_state[10] <<< 0;
wire signed [31:0] shifted_state198_10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state198_10_2 = reservoir_state[10] <<< 2;
wire signed [31:0] shifted_state198_10_3 = reservoir_state[10] <<< 3;
wire signed [31:0] shifted_state198_10_4 = reservoir_state[10] <<< 4;
wire signed [31:0] shifted_state198_10_5 = reservoir_state[10] <<< 5;
wire signed [31:0] shifted_state198_10_6 = reservoir_state[10] <<< 6;
wire signed [31:0] shifted_state198_10_7 = reservoir_state[10] <<< 7;
wire signed [31:0] shifted_state198_11_1 = reservoir_state[11] <<< 1;
wire signed [31:0] shifted_state198_11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state198_11_3 = reservoir_state[11] <<< 3;
wire signed [31:0] shifted_state198_11_4 = reservoir_state[11] <<< 4;
wire signed [31:0] shifted_state198_24_0 = reservoir_state[24] <<< 0;
wire signed [31:0] shifted_state198_24_2 = reservoir_state[24] <<< 2;
wire signed [31:0] shifted_state198_24_4 = reservoir_state[24] <<< 4;
wire signed [31:0] shifted_state198_42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state198_42_2 = reservoir_state[42] <<< 2;
wire signed [31:0] shifted_state198_42_4 = reservoir_state[42] <<< 4;
wire signed [31:0] shifted_state198_83_1 = reservoir_state[83] <<< 1;
wire signed [31:0] shifted_state198_83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state198_83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state198_83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state198_83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state198_84_0 = reservoir_state[84] <<< 0;
wire signed [31:0] shifted_state198_84_1 = reservoir_state[84] <<< 1;
wire signed [31:0] shifted_state198_84_5 = reservoir_state[84] <<< 5;
wire signed [31:0] shifted_state198_84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state198_84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state198_105_3 = reservoir_state[105] <<< 3;
wire signed [31:0] shifted_state198_105_4 = reservoir_state[105] <<< 4;
wire signed [31:0] shifted_state198_105_5 = reservoir_state[105] <<< 5;
wire signed [31:0] shifted_state198_105_6 = reservoir_state[105] <<< 6;
wire signed [31:0] shifted_state198_105_7 = reservoir_state[105] <<< 7;
wire signed [31:0] shifted_state198_116_1 = reservoir_state[116] <<< 1;
wire signed [31:0] shifted_state198_116_2 = reservoir_state[116] <<< 2;
wire signed [31:0] shifted_state198_116_3 = reservoir_state[116] <<< 3;
wire signed [31:0] shifted_state198_116_4 = reservoir_state[116] <<< 4;
wire signed [31:0] shifted_state198_116_5 = reservoir_state[116] <<< 5;
wire signed [31:0] shifted_state198_116_6 = reservoir_state[116] <<< 6;
wire signed [31:0] shifted_state198_116_7 = reservoir_state[116] <<< 7;
wire signed [31:0] shifted_state198_128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state198_152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state198_152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state198_158_1 = reservoir_state[158] <<< 1;
wire signed [31:0] shifted_state198_158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state198_158_3 = reservoir_state[158] <<< 3;
wire signed [31:0] shifted_state198_158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state198_158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state198_158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state198_158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state198_160_1 = reservoir_state[160] <<< 1;
wire signed [31:0] shifted_state198_160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state198_160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state198_160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state198_160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state198_161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state198_161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state198_161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state198_161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state198_161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state198_161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state198_179_0 = reservoir_state[179] <<< 0;
wire signed [31:0] shifted_state198_179_1 = reservoir_state[179] <<< 1;
wire signed [31:0] shifted_state198_179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state198_179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state198_179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state198_179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state198_188_1 = reservoir_state[188] <<< 1;
wire signed [31:0] shifted_state198_188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state198_188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state198_188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state198_188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state198_188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state198_188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state198_189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state198_189_2 = reservoir_state[189] <<< 2;
wire signed [31:0] shifted_state198_189_3 = reservoir_state[189] <<< 3;
wire signed [31:0] shifted_state198_189_4 = reservoir_state[189] <<< 4;
wire signed [31:0] shifted_state199_2_1 = reservoir_state[2] <<< 1;
wire signed [31:0] shifted_state199_2_4 = reservoir_state[2] <<< 4;
wire signed [31:0] shifted_state199_6_0 = reservoir_state[6] <<< 0;
wire signed [31:0] shifted_state199_6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state199_6_2 = reservoir_state[6] <<< 2;
wire signed [31:0] shifted_state199_6_5 = reservoir_state[6] <<< 5;
wire signed [31:0] shifted_state199_41_0 = reservoir_state[41] <<< 0;
wire signed [31:0] shifted_state199_41_2 = reservoir_state[41] <<< 2;
wire signed [31:0] shifted_state199_41_4 = reservoir_state[41] <<< 4;
wire signed [31:0] shifted_state199_41_6 = reservoir_state[41] <<< 6;
wire signed [31:0] shifted_state199_41_7 = reservoir_state[41] <<< 7;
wire signed [31:0] shifted_state199_53_1 = reservoir_state[53] <<< 1;
wire signed [31:0] shifted_state199_53_3 = reservoir_state[53] <<< 3;
wire signed [31:0] shifted_state199_59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state199_59_2 = reservoir_state[59] <<< 2;
wire signed [31:0] shifted_state199_59_4 = reservoir_state[59] <<< 4;
wire signed [31:0] shifted_state199_59_6 = reservoir_state[59] <<< 6;
wire signed [31:0] shifted_state199_59_7 = reservoir_state[59] <<< 7;
wire signed [31:0] shifted_state199_64_0 = reservoir_state[64] <<< 0;
wire signed [31:0] shifted_state199_64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state199_65_1 = reservoir_state[65] <<< 1;
wire signed [31:0] shifted_state199_65_2 = reservoir_state[65] <<< 2;
wire signed [31:0] shifted_state199_65_4 = reservoir_state[65] <<< 4;
wire signed [31:0] shifted_state199_78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state199_82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state199_82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state199_82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state199_82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state199_136_0 = reservoir_state[136] <<< 0;
wire signed [31:0] shifted_state199_136_4 = reservoir_state[136] <<< 4;
wire signed [31:0] shifted_state199_136_5 = reservoir_state[136] <<< 5;
wire signed [31:0] shifted_state199_145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state199_145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state199_145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state199_145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state199_145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state199_146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state199_146_2 = reservoir_state[146] <<< 2;
wire signed [31:0] shifted_state199_146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state199_159_2 = reservoir_state[159] <<< 2;
wire signed [31:0] shifted_state199_159_3 = reservoir_state[159] <<< 3;
wire signed [31:0] shifted_state199_159_4 = reservoir_state[159] <<< 4;
wire signed [31:0] shifted_state199_159_5 = reservoir_state[159] <<< 5;
wire signed [31:0] shifted_state199_159_6 = reservoir_state[159] <<< 6;
wire signed [31:0] shifted_state199_159_7 = reservoir_state[159] <<< 7;
wire signed [31:0] shifted_state199_176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state199_176_2 = reservoir_state[176] <<< 2;
wire signed [31:0] shifted_state199_176_4 = reservoir_state[176] <<< 4;
wire signed [31:0] shifted_state199_186_1 = reservoir_state[186] <<< 1;
wire signed [31:0] shifted_state199_186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state199_186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state199_186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state199_186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state199_186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state199_186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state199_191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state199_191_5 = reservoir_state[191] <<< 5;
wire signed [31:0] shifted_state199_191_6 = reservoir_state[191] <<< 6;
wire signed [31:0] shifted_state199_191_7 = reservoir_state[191] <<< 7;
wire signed [31:0] shifted_state_out0_0 = reservoir_state[0] <<< 0;
wire signed [31:0] shifted_state_out0_2 = reservoir_state[0] <<< 2;
wire signed [31:0] shifted_state_out0_3 = reservoir_state[0] <<< 3;
wire signed [31:0] shifted_state_out0_4 = reservoir_state[0] <<< 4;
wire signed [31:0] shifted_state_out0_5 = reservoir_state[0] <<< 5;
wire signed [31:0] shifted_state_out0_6 = reservoir_state[0] <<< 6;
wire signed [31:0] shifted_state_out0_7 = reservoir_state[0] <<< 7;
wire signed [31:0] shifted_state_out1_0 = reservoir_state[1] <<< 0;
wire signed [31:0] shifted_state_out1_2 = reservoir_state[1] <<< 2;
wire signed [31:0] shifted_state_out2_2 = reservoir_state[2] <<< 2;
wire signed [31:0] shifted_state_out3_1 = reservoir_state[3] <<< 1;
wire signed [31:0] shifted_state_out5_1 = reservoir_state[5] <<< 1;
wire signed [31:0] shifted_state_out5_2 = reservoir_state[5] <<< 2;
wire signed [31:0] shifted_state_out5_3 = reservoir_state[5] <<< 3;
wire signed [31:0] shifted_state_out5_4 = reservoir_state[5] <<< 4;
wire signed [31:0] shifted_state_out5_5 = reservoir_state[5] <<< 5;
wire signed [31:0] shifted_state_out5_6 = reservoir_state[5] <<< 6;
wire signed [31:0] shifted_state_out5_7 = reservoir_state[5] <<< 7;
wire signed [31:0] shifted_state_out6_1 = reservoir_state[6] <<< 1;
wire signed [31:0] shifted_state_out7_1 = reservoir_state[7] <<< 1;
wire signed [31:0] shifted_state_out7_3 = reservoir_state[7] <<< 3;
wire signed [31:0] shifted_state_out7_4 = reservoir_state[7] <<< 4;
wire signed [31:0] shifted_state_out7_5 = reservoir_state[7] <<< 5;
wire signed [31:0] shifted_state_out7_6 = reservoir_state[7] <<< 6;
wire signed [31:0] shifted_state_out7_7 = reservoir_state[7] <<< 7;
wire signed [31:0] shifted_state_out9_2 = reservoir_state[9] <<< 2;
wire signed [31:0] shifted_state_out10_1 = reservoir_state[10] <<< 1;
wire signed [31:0] shifted_state_out11_0 = reservoir_state[11] <<< 0;
wire signed [31:0] shifted_state_out11_2 = reservoir_state[11] <<< 2;
wire signed [31:0] shifted_state_out12_1 = reservoir_state[12] <<< 1;
wire signed [31:0] shifted_state_out13_0 = reservoir_state[13] <<< 0;
wire signed [31:0] shifted_state_out13_2 = reservoir_state[13] <<< 2;
wire signed [31:0] shifted_state_out13_3 = reservoir_state[13] <<< 3;
wire signed [31:0] shifted_state_out13_4 = reservoir_state[13] <<< 4;
wire signed [31:0] shifted_state_out13_5 = reservoir_state[13] <<< 5;
wire signed [31:0] shifted_state_out13_6 = reservoir_state[13] <<< 6;
wire signed [31:0] shifted_state_out13_7 = reservoir_state[13] <<< 7;
wire signed [31:0] shifted_state_out14_0 = reservoir_state[14] <<< 0;
wire signed [31:0] shifted_state_out14_1 = reservoir_state[14] <<< 1;
wire signed [31:0] shifted_state_out15_0 = reservoir_state[15] <<< 0;
wire signed [31:0] shifted_state_out15_4 = reservoir_state[15] <<< 4;
wire signed [31:0] shifted_state_out16_0 = reservoir_state[16] <<< 0;
wire signed [31:0] shifted_state_out16_2 = reservoir_state[16] <<< 2;
wire signed [31:0] shifted_state_out16_4 = reservoir_state[16] <<< 4;
wire signed [31:0] shifted_state_out16_5 = reservoir_state[16] <<< 5;
wire signed [31:0] shifted_state_out16_6 = reservoir_state[16] <<< 6;
wire signed [31:0] shifted_state_out16_7 = reservoir_state[16] <<< 7;
wire signed [31:0] shifted_state_out17_1 = reservoir_state[17] <<< 1;
wire signed [31:0] shifted_state_out17_2 = reservoir_state[17] <<< 2;
wire signed [31:0] shifted_state_out17_3 = reservoir_state[17] <<< 3;
wire signed [31:0] shifted_state_out17_4 = reservoir_state[17] <<< 4;
wire signed [31:0] shifted_state_out17_5 = reservoir_state[17] <<< 5;
wire signed [31:0] shifted_state_out17_6 = reservoir_state[17] <<< 6;
wire signed [31:0] shifted_state_out17_7 = reservoir_state[17] <<< 7;
wire signed [31:0] shifted_state_out18_0 = reservoir_state[18] <<< 0;
wire signed [31:0] shifted_state_out18_1 = reservoir_state[18] <<< 1;
wire signed [31:0] shifted_state_out19_0 = reservoir_state[19] <<< 0;
wire signed [31:0] shifted_state_out19_1 = reservoir_state[19] <<< 1;
wire signed [31:0] shifted_state_out19_2 = reservoir_state[19] <<< 2;
wire signed [31:0] shifted_state_out19_3 = reservoir_state[19] <<< 3;
wire signed [31:0] shifted_state_out20_2 = reservoir_state[20] <<< 2;
wire signed [31:0] shifted_state_out21_0 = reservoir_state[21] <<< 0;
wire signed [31:0] shifted_state_out21_1 = reservoir_state[21] <<< 1;
wire signed [31:0] shifted_state_out21_2 = reservoir_state[21] <<< 2;
wire signed [31:0] shifted_state_out21_3 = reservoir_state[21] <<< 3;
wire signed [31:0] shifted_state_out21_4 = reservoir_state[21] <<< 4;
wire signed [31:0] shifted_state_out21_5 = reservoir_state[21] <<< 5;
wire signed [31:0] shifted_state_out21_6 = reservoir_state[21] <<< 6;
wire signed [31:0] shifted_state_out21_7 = reservoir_state[21] <<< 7;
wire signed [31:0] shifted_state_out22_0 = reservoir_state[22] <<< 0;
wire signed [31:0] shifted_state_out22_1 = reservoir_state[22] <<< 1;
wire signed [31:0] shifted_state_out23_3 = reservoir_state[23] <<< 3;
wire signed [31:0] shifted_state_out24_1 = reservoir_state[24] <<< 1;
wire signed [31:0] shifted_state_out25_1 = reservoir_state[25] <<< 1;
wire signed [31:0] shifted_state_out25_4 = reservoir_state[25] <<< 4;
wire signed [31:0] shifted_state_out25_5 = reservoir_state[25] <<< 5;
wire signed [31:0] shifted_state_out26_1 = reservoir_state[26] <<< 1;
wire signed [31:0] shifted_state_out26_2 = reservoir_state[26] <<< 2;
wire signed [31:0] shifted_state_out27_1 = reservoir_state[27] <<< 1;
wire signed [31:0] shifted_state_out27_2 = reservoir_state[27] <<< 2;
wire signed [31:0] shifted_state_out28_0 = reservoir_state[28] <<< 0;
wire signed [31:0] shifted_state_out28_2 = reservoir_state[28] <<< 2;
wire signed [31:0] shifted_state_out30_1 = reservoir_state[30] <<< 1;
wire signed [31:0] shifted_state_out30_2 = reservoir_state[30] <<< 2;
wire signed [31:0] shifted_state_out30_3 = reservoir_state[30] <<< 3;
wire signed [31:0] shifted_state_out30_4 = reservoir_state[30] <<< 4;
wire signed [31:0] shifted_state_out30_5 = reservoir_state[30] <<< 5;
wire signed [31:0] shifted_state_out30_6 = reservoir_state[30] <<< 6;
wire signed [31:0] shifted_state_out30_7 = reservoir_state[30] <<< 7;
wire signed [31:0] shifted_state_out31_3 = reservoir_state[31] <<< 3;
wire signed [31:0] shifted_state_out32_0 = reservoir_state[32] <<< 0;
wire signed [31:0] shifted_state_out32_1 = reservoir_state[32] <<< 1;
wire signed [31:0] shifted_state_out32_3 = reservoir_state[32] <<< 3;
wire signed [31:0] shifted_state_out32_4 = reservoir_state[32] <<< 4;
wire signed [31:0] shifted_state_out32_5 = reservoir_state[32] <<< 5;
wire signed [31:0] shifted_state_out32_6 = reservoir_state[32] <<< 6;
wire signed [31:0] shifted_state_out32_7 = reservoir_state[32] <<< 7;
wire signed [31:0] shifted_state_out33_1 = reservoir_state[33] <<< 1;
wire signed [31:0] shifted_state_out34_2 = reservoir_state[34] <<< 2;
wire signed [31:0] shifted_state_out35_0 = reservoir_state[35] <<< 0;
wire signed [31:0] shifted_state_out35_1 = reservoir_state[35] <<< 1;
wire signed [31:0] shifted_state_out35_2 = reservoir_state[35] <<< 2;
wire signed [31:0] shifted_state_out36_1 = reservoir_state[36] <<< 1;
wire signed [31:0] shifted_state_out36_2 = reservoir_state[36] <<< 2;
wire signed [31:0] shifted_state_out36_3 = reservoir_state[36] <<< 3;
wire signed [31:0] shifted_state_out36_4 = reservoir_state[36] <<< 4;
wire signed [31:0] shifted_state_out36_5 = reservoir_state[36] <<< 5;
wire signed [31:0] shifted_state_out36_6 = reservoir_state[36] <<< 6;
wire signed [31:0] shifted_state_out36_7 = reservoir_state[36] <<< 7;
wire signed [31:0] shifted_state_out37_0 = reservoir_state[37] <<< 0;
wire signed [31:0] shifted_state_out37_1 = reservoir_state[37] <<< 1;
wire signed [31:0] shifted_state_out38_1 = reservoir_state[38] <<< 1;
wire signed [31:0] shifted_state_out38_3 = reservoir_state[38] <<< 3;
wire signed [31:0] shifted_state_out38_4 = reservoir_state[38] <<< 4;
wire signed [31:0] shifted_state_out38_5 = reservoir_state[38] <<< 5;
wire signed [31:0] shifted_state_out38_6 = reservoir_state[38] <<< 6;
wire signed [31:0] shifted_state_out38_7 = reservoir_state[38] <<< 7;
wire signed [31:0] shifted_state_out39_1 = reservoir_state[39] <<< 1;
wire signed [31:0] shifted_state_out39_3 = reservoir_state[39] <<< 3;
wire signed [31:0] shifted_state_out39_4 = reservoir_state[39] <<< 4;
wire signed [31:0] shifted_state_out39_5 = reservoir_state[39] <<< 5;
wire signed [31:0] shifted_state_out39_6 = reservoir_state[39] <<< 6;
wire signed [31:0] shifted_state_out39_7 = reservoir_state[39] <<< 7;
wire signed [31:0] shifted_state_out40_1 = reservoir_state[40] <<< 1;
wire signed [31:0] shifted_state_out42_0 = reservoir_state[42] <<< 0;
wire signed [31:0] shifted_state_out42_3 = reservoir_state[42] <<< 3;
wire signed [31:0] shifted_state_out43_0 = reservoir_state[43] <<< 0;
wire signed [31:0] shifted_state_out43_1 = reservoir_state[43] <<< 1;
wire signed [31:0] shifted_state_out43_2 = reservoir_state[43] <<< 2;
wire signed [31:0] shifted_state_out43_3 = reservoir_state[43] <<< 3;
wire signed [31:0] shifted_state_out43_4 = reservoir_state[43] <<< 4;
wire signed [31:0] shifted_state_out43_5 = reservoir_state[43] <<< 5;
wire signed [31:0] shifted_state_out43_6 = reservoir_state[43] <<< 6;
wire signed [31:0] shifted_state_out43_7 = reservoir_state[43] <<< 7;
wire signed [31:0] shifted_state_out44_1 = reservoir_state[44] <<< 1;
wire signed [31:0] shifted_state_out45_2 = reservoir_state[45] <<< 2;
wire signed [31:0] shifted_state_out45_3 = reservoir_state[45] <<< 3;
wire signed [31:0] shifted_state_out45_4 = reservoir_state[45] <<< 4;
wire signed [31:0] shifted_state_out45_5 = reservoir_state[45] <<< 5;
wire signed [31:0] shifted_state_out45_6 = reservoir_state[45] <<< 6;
wire signed [31:0] shifted_state_out45_7 = reservoir_state[45] <<< 7;
wire signed [31:0] shifted_state_out46_0 = reservoir_state[46] <<< 0;
wire signed [31:0] shifted_state_out46_3 = reservoir_state[46] <<< 3;
wire signed [31:0] shifted_state_out46_4 = reservoir_state[46] <<< 4;
wire signed [31:0] shifted_state_out46_5 = reservoir_state[46] <<< 5;
wire signed [31:0] shifted_state_out46_6 = reservoir_state[46] <<< 6;
wire signed [31:0] shifted_state_out46_7 = reservoir_state[46] <<< 7;
wire signed [31:0] shifted_state_out47_0 = reservoir_state[47] <<< 0;
wire signed [31:0] shifted_state_out47_1 = reservoir_state[47] <<< 1;
wire signed [31:0] shifted_state_out48_1 = reservoir_state[48] <<< 1;
wire signed [31:0] shifted_state_out48_2 = reservoir_state[48] <<< 2;
wire signed [31:0] shifted_state_out48_3 = reservoir_state[48] <<< 3;
wire signed [31:0] shifted_state_out48_4 = reservoir_state[48] <<< 4;
wire signed [31:0] shifted_state_out48_5 = reservoir_state[48] <<< 5;
wire signed [31:0] shifted_state_out48_6 = reservoir_state[48] <<< 6;
wire signed [31:0] shifted_state_out48_7 = reservoir_state[48] <<< 7;
wire signed [31:0] shifted_state_out50_1 = reservoir_state[50] <<< 1;
wire signed [31:0] shifted_state_out50_2 = reservoir_state[50] <<< 2;
wire signed [31:0] shifted_state_out51_0 = reservoir_state[51] <<< 0;
wire signed [31:0] shifted_state_out51_3 = reservoir_state[51] <<< 3;
wire signed [31:0] shifted_state_out52_0 = reservoir_state[52] <<< 0;
wire signed [31:0] shifted_state_out52_2 = reservoir_state[52] <<< 2;
wire signed [31:0] shifted_state_out52_3 = reservoir_state[52] <<< 3;
wire signed [31:0] shifted_state_out52_4 = reservoir_state[52] <<< 4;
wire signed [31:0] shifted_state_out52_5 = reservoir_state[52] <<< 5;
wire signed [31:0] shifted_state_out52_6 = reservoir_state[52] <<< 6;
wire signed [31:0] shifted_state_out52_7 = reservoir_state[52] <<< 7;
wire signed [31:0] shifted_state_out53_0 = reservoir_state[53] <<< 0;
wire signed [31:0] shifted_state_out53_1 = reservoir_state[53] <<< 1;
wire signed [31:0] shifted_state_out53_2 = reservoir_state[53] <<< 2;
wire signed [31:0] shifted_state_out55_0 = reservoir_state[55] <<< 0;
wire signed [31:0] shifted_state_out55_1 = reservoir_state[55] <<< 1;
wire signed [31:0] shifted_state_out55_3 = reservoir_state[55] <<< 3;
wire signed [31:0] shifted_state_out55_4 = reservoir_state[55] <<< 4;
wire signed [31:0] shifted_state_out55_5 = reservoir_state[55] <<< 5;
wire signed [31:0] shifted_state_out55_6 = reservoir_state[55] <<< 6;
wire signed [31:0] shifted_state_out55_7 = reservoir_state[55] <<< 7;
wire signed [31:0] shifted_state_out56_1 = reservoir_state[56] <<< 1;
wire signed [31:0] shifted_state_out57_0 = reservoir_state[57] <<< 0;
wire signed [31:0] shifted_state_out57_1 = reservoir_state[57] <<< 1;
wire signed [31:0] shifted_state_out57_2 = reservoir_state[57] <<< 2;
wire signed [31:0] shifted_state_out58_0 = reservoir_state[58] <<< 0;
wire signed [31:0] shifted_state_out58_2 = reservoir_state[58] <<< 2;
wire signed [31:0] shifted_state_out58_3 = reservoir_state[58] <<< 3;
wire signed [31:0] shifted_state_out58_4 = reservoir_state[58] <<< 4;
wire signed [31:0] shifted_state_out58_5 = reservoir_state[58] <<< 5;
wire signed [31:0] shifted_state_out58_6 = reservoir_state[58] <<< 6;
wire signed [31:0] shifted_state_out58_7 = reservoir_state[58] <<< 7;
wire signed [31:0] shifted_state_out59_0 = reservoir_state[59] <<< 0;
wire signed [31:0] shifted_state_out59_1 = reservoir_state[59] <<< 1;
wire signed [31:0] shifted_state_out61_0 = reservoir_state[61] <<< 0;
wire signed [31:0] shifted_state_out62_1 = reservoir_state[62] <<< 1;
wire signed [31:0] shifted_state_out62_2 = reservoir_state[62] <<< 2;
wire signed [31:0] shifted_state_out62_3 = reservoir_state[62] <<< 3;
wire signed [31:0] shifted_state_out62_4 = reservoir_state[62] <<< 4;
wire signed [31:0] shifted_state_out62_5 = reservoir_state[62] <<< 5;
wire signed [31:0] shifted_state_out62_6 = reservoir_state[62] <<< 6;
wire signed [31:0] shifted_state_out62_7 = reservoir_state[62] <<< 7;
wire signed [31:0] shifted_state_out63_3 = reservoir_state[63] <<< 3;
wire signed [31:0] shifted_state_out64_1 = reservoir_state[64] <<< 1;
wire signed [31:0] shifted_state_out64_2 = reservoir_state[64] <<< 2;
wire signed [31:0] shifted_state_out64_3 = reservoir_state[64] <<< 3;
wire signed [31:0] shifted_state_out64_4 = reservoir_state[64] <<< 4;
wire signed [31:0] shifted_state_out64_5 = reservoir_state[64] <<< 5;
wire signed [31:0] shifted_state_out64_6 = reservoir_state[64] <<< 6;
wire signed [31:0] shifted_state_out64_7 = reservoir_state[64] <<< 7;
wire signed [31:0] shifted_state_out65_0 = reservoir_state[65] <<< 0;
wire signed [31:0] shifted_state_out65_2 = reservoir_state[65] <<< 2;
wire signed [31:0] shifted_state_out66_1 = reservoir_state[66] <<< 1;
wire signed [31:0] shifted_state_out67_0 = reservoir_state[67] <<< 0;
wire signed [31:0] shifted_state_out69_0 = reservoir_state[69] <<< 0;
wire signed [31:0] shifted_state_out70_1 = reservoir_state[70] <<< 1;
wire signed [31:0] shifted_state_out70_3 = reservoir_state[70] <<< 3;
wire signed [31:0] shifted_state_out70_4 = reservoir_state[70] <<< 4;
wire signed [31:0] shifted_state_out70_5 = reservoir_state[70] <<< 5;
wire signed [31:0] shifted_state_out70_6 = reservoir_state[70] <<< 6;
wire signed [31:0] shifted_state_out70_7 = reservoir_state[70] <<< 7;
wire signed [31:0] shifted_state_out71_1 = reservoir_state[71] <<< 1;
wire signed [31:0] shifted_state_out72_0 = reservoir_state[72] <<< 0;
wire signed [31:0] shifted_state_out72_1 = reservoir_state[72] <<< 1;
wire signed [31:0] shifted_state_out72_3 = reservoir_state[72] <<< 3;
wire signed [31:0] shifted_state_out72_4 = reservoir_state[72] <<< 4;
wire signed [31:0] shifted_state_out72_5 = reservoir_state[72] <<< 5;
wire signed [31:0] shifted_state_out72_6 = reservoir_state[72] <<< 6;
wire signed [31:0] shifted_state_out72_7 = reservoir_state[72] <<< 7;
wire signed [31:0] shifted_state_out73_0 = reservoir_state[73] <<< 0;
wire signed [31:0] shifted_state_out73_1 = reservoir_state[73] <<< 1;
wire signed [31:0] shifted_state_out73_3 = reservoir_state[73] <<< 3;
wire signed [31:0] shifted_state_out73_4 = reservoir_state[73] <<< 4;
wire signed [31:0] shifted_state_out73_5 = reservoir_state[73] <<< 5;
wire signed [31:0] shifted_state_out73_6 = reservoir_state[73] <<< 6;
wire signed [31:0] shifted_state_out73_7 = reservoir_state[73] <<< 7;
wire signed [31:0] shifted_state_out74_0 = reservoir_state[74] <<< 0;
wire signed [31:0] shifted_state_out74_2 = reservoir_state[74] <<< 2;
wire signed [31:0] shifted_state_out75_0 = reservoir_state[75] <<< 0;
wire signed [31:0] shifted_state_out76_1 = reservoir_state[76] <<< 1;
wire signed [31:0] shifted_state_out76_2 = reservoir_state[76] <<< 2;
wire signed [31:0] shifted_state_out76_3 = reservoir_state[76] <<< 3;
wire signed [31:0] shifted_state_out76_4 = reservoir_state[76] <<< 4;
wire signed [31:0] shifted_state_out76_5 = reservoir_state[76] <<< 5;
wire signed [31:0] shifted_state_out76_6 = reservoir_state[76] <<< 6;
wire signed [31:0] shifted_state_out76_7 = reservoir_state[76] <<< 7;
wire signed [31:0] shifted_state_out77_2 = reservoir_state[77] <<< 2;
wire signed [31:0] shifted_state_out77_3 = reservoir_state[77] <<< 3;
wire signed [31:0] shifted_state_out77_4 = reservoir_state[77] <<< 4;
wire signed [31:0] shifted_state_out77_5 = reservoir_state[77] <<< 5;
wire signed [31:0] shifted_state_out77_6 = reservoir_state[77] <<< 6;
wire signed [31:0] shifted_state_out77_7 = reservoir_state[77] <<< 7;
wire signed [31:0] shifted_state_out78_0 = reservoir_state[78] <<< 0;
wire signed [31:0] shifted_state_out78_1 = reservoir_state[78] <<< 1;
wire signed [31:0] shifted_state_out78_2 = reservoir_state[78] <<< 2;
wire signed [31:0] shifted_state_out78_3 = reservoir_state[78] <<< 3;
wire signed [31:0] shifted_state_out78_4 = reservoir_state[78] <<< 4;
wire signed [31:0] shifted_state_out78_5 = reservoir_state[78] <<< 5;
wire signed [31:0] shifted_state_out78_6 = reservoir_state[78] <<< 6;
wire signed [31:0] shifted_state_out78_7 = reservoir_state[78] <<< 7;
wire signed [31:0] shifted_state_out79_1 = reservoir_state[79] <<< 1;
wire signed [31:0] shifted_state_out79_2 = reservoir_state[79] <<< 2;
wire signed [31:0] shifted_state_out79_3 = reservoir_state[79] <<< 3;
wire signed [31:0] shifted_state_out79_4 = reservoir_state[79] <<< 4;
wire signed [31:0] shifted_state_out79_5 = reservoir_state[79] <<< 5;
wire signed [31:0] shifted_state_out79_6 = reservoir_state[79] <<< 6;
wire signed [31:0] shifted_state_out79_7 = reservoir_state[79] <<< 7;
wire signed [31:0] shifted_state_out80_0 = reservoir_state[80] <<< 0;
wire signed [31:0] shifted_state_out80_1 = reservoir_state[80] <<< 1;
wire signed [31:0] shifted_state_out80_2 = reservoir_state[80] <<< 2;
wire signed [31:0] shifted_state_out81_0 = reservoir_state[81] <<< 0;
wire signed [31:0] shifted_state_out82_0 = reservoir_state[82] <<< 0;
wire signed [31:0] shifted_state_out82_1 = reservoir_state[82] <<< 1;
wire signed [31:0] shifted_state_out82_2 = reservoir_state[82] <<< 2;
wire signed [31:0] shifted_state_out82_3 = reservoir_state[82] <<< 3;
wire signed [31:0] shifted_state_out82_4 = reservoir_state[82] <<< 4;
wire signed [31:0] shifted_state_out82_5 = reservoir_state[82] <<< 5;
wire signed [31:0] shifted_state_out82_6 = reservoir_state[82] <<< 6;
wire signed [31:0] shifted_state_out82_7 = reservoir_state[82] <<< 7;
wire signed [31:0] shifted_state_out83_2 = reservoir_state[83] <<< 2;
wire signed [31:0] shifted_state_out83_3 = reservoir_state[83] <<< 3;
wire signed [31:0] shifted_state_out83_4 = reservoir_state[83] <<< 4;
wire signed [31:0] shifted_state_out83_5 = reservoir_state[83] <<< 5;
wire signed [31:0] shifted_state_out83_6 = reservoir_state[83] <<< 6;
wire signed [31:0] shifted_state_out83_7 = reservoir_state[83] <<< 7;
wire signed [31:0] shifted_state_out84_3 = reservoir_state[84] <<< 3;
wire signed [31:0] shifted_state_out84_4 = reservoir_state[84] <<< 4;
wire signed [31:0] shifted_state_out84_5 = reservoir_state[84] <<< 5;
wire signed [31:0] shifted_state_out84_6 = reservoir_state[84] <<< 6;
wire signed [31:0] shifted_state_out84_7 = reservoir_state[84] <<< 7;
wire signed [31:0] shifted_state_out85_0 = reservoir_state[85] <<< 0;
wire signed [31:0] shifted_state_out86_2 = reservoir_state[86] <<< 2;
wire signed [31:0] shifted_state_out87_3 = reservoir_state[87] <<< 3;
wire signed [31:0] shifted_state_out87_4 = reservoir_state[87] <<< 4;
wire signed [31:0] shifted_state_out87_5 = reservoir_state[87] <<< 5;
wire signed [31:0] shifted_state_out87_6 = reservoir_state[87] <<< 6;
wire signed [31:0] shifted_state_out87_7 = reservoir_state[87] <<< 7;
wire signed [31:0] shifted_state_out88_0 = reservoir_state[88] <<< 0;
wire signed [31:0] shifted_state_out89_2 = reservoir_state[89] <<< 2;
wire signed [31:0] shifted_state_out89_3 = reservoir_state[89] <<< 3;
wire signed [31:0] shifted_state_out90_3 = reservoir_state[90] <<< 3;
wire signed [31:0] shifted_state_out91_0 = reservoir_state[91] <<< 0;
wire signed [31:0] shifted_state_out91_1 = reservoir_state[91] <<< 1;
wire signed [31:0] shifted_state_out91_3 = reservoir_state[91] <<< 3;
wire signed [31:0] shifted_state_out91_4 = reservoir_state[91] <<< 4;
wire signed [31:0] shifted_state_out91_5 = reservoir_state[91] <<< 5;
wire signed [31:0] shifted_state_out91_6 = reservoir_state[91] <<< 6;
wire signed [31:0] shifted_state_out91_7 = reservoir_state[91] <<< 7;
wire signed [31:0] shifted_state_out92_0 = reservoir_state[92] <<< 0;
wire signed [31:0] shifted_state_out92_2 = reservoir_state[92] <<< 2;
wire signed [31:0] shifted_state_out93_0 = reservoir_state[93] <<< 0;
wire signed [31:0] shifted_state_out93_1 = reservoir_state[93] <<< 1;
wire signed [31:0] shifted_state_out93_2 = reservoir_state[93] <<< 2;
wire signed [31:0] shifted_state_out93_3 = reservoir_state[93] <<< 3;
wire signed [31:0] shifted_state_out93_4 = reservoir_state[93] <<< 4;
wire signed [31:0] shifted_state_out93_5 = reservoir_state[93] <<< 5;
wire signed [31:0] shifted_state_out93_6 = reservoir_state[93] <<< 6;
wire signed [31:0] shifted_state_out93_7 = reservoir_state[93] <<< 7;
wire signed [31:0] shifted_state_out95_0 = reservoir_state[95] <<< 0;
wire signed [31:0] shifted_state_out95_1 = reservoir_state[95] <<< 1;
wire signed [31:0] shifted_state_out95_2 = reservoir_state[95] <<< 2;
wire signed [31:0] shifted_state_out95_3 = reservoir_state[95] <<< 3;
wire signed [31:0] shifted_state_out95_4 = reservoir_state[95] <<< 4;
wire signed [31:0] shifted_state_out95_5 = reservoir_state[95] <<< 5;
wire signed [31:0] shifted_state_out95_6 = reservoir_state[95] <<< 6;
wire signed [31:0] shifted_state_out95_7 = reservoir_state[95] <<< 7;
wire signed [31:0] shifted_state_out96_0 = reservoir_state[96] <<< 0;
wire signed [31:0] shifted_state_out96_2 = reservoir_state[96] <<< 2;
wire signed [31:0] shifted_state_out97_0 = reservoir_state[97] <<< 0;
wire signed [31:0] shifted_state_out97_1 = reservoir_state[97] <<< 1;
wire signed [31:0] shifted_state_out97_2 = reservoir_state[97] <<< 2;
wire signed [31:0] shifted_state_out97_3 = reservoir_state[97] <<< 3;
wire signed [31:0] shifted_state_out97_4 = reservoir_state[97] <<< 4;
wire signed [31:0] shifted_state_out97_5 = reservoir_state[97] <<< 5;
wire signed [31:0] shifted_state_out97_6 = reservoir_state[97] <<< 6;
wire signed [31:0] shifted_state_out97_7 = reservoir_state[97] <<< 7;
wire signed [31:0] shifted_state_out98_2 = reservoir_state[98] <<< 2;
wire signed [31:0] shifted_state_out100_0 = reservoir_state[100] <<< 0;
wire signed [31:0] shifted_state_out100_1 = reservoir_state[100] <<< 1;
wire signed [31:0] shifted_state_out100_3 = reservoir_state[100] <<< 3;
wire signed [31:0] shifted_state_out100_4 = reservoir_state[100] <<< 4;
wire signed [31:0] shifted_state_out100_5 = reservoir_state[100] <<< 5;
wire signed [31:0] shifted_state_out100_6 = reservoir_state[100] <<< 6;
wire signed [31:0] shifted_state_out100_7 = reservoir_state[100] <<< 7;
wire signed [31:0] shifted_state_out101_1 = reservoir_state[101] <<< 1;
wire signed [31:0] shifted_state_out102_1 = reservoir_state[102] <<< 1;
wire signed [31:0] shifted_state_out102_2 = reservoir_state[102] <<< 2;
wire signed [31:0] shifted_state_out102_3 = reservoir_state[102] <<< 3;
wire signed [31:0] shifted_state_out102_4 = reservoir_state[102] <<< 4;
wire signed [31:0] shifted_state_out102_5 = reservoir_state[102] <<< 5;
wire signed [31:0] shifted_state_out102_6 = reservoir_state[102] <<< 6;
wire signed [31:0] shifted_state_out102_7 = reservoir_state[102] <<< 7;
wire signed [31:0] shifted_state_out103_1 = reservoir_state[103] <<< 1;
wire signed [31:0] shifted_state_out103_2 = reservoir_state[103] <<< 2;
wire signed [31:0] shifted_state_out103_3 = reservoir_state[103] <<< 3;
wire signed [31:0] shifted_state_out103_4 = reservoir_state[103] <<< 4;
wire signed [31:0] shifted_state_out103_5 = reservoir_state[103] <<< 5;
wire signed [31:0] shifted_state_out103_6 = reservoir_state[103] <<< 6;
wire signed [31:0] shifted_state_out103_7 = reservoir_state[103] <<< 7;
wire signed [31:0] shifted_state_out105_0 = reservoir_state[105] <<< 0;
wire signed [31:0] shifted_state_out105_2 = reservoir_state[105] <<< 2;
wire signed [31:0] shifted_state_out106_0 = reservoir_state[106] <<< 0;
wire signed [31:0] shifted_state_out106_1 = reservoir_state[106] <<< 1;
wire signed [31:0] shifted_state_out107_0 = reservoir_state[107] <<< 0;
wire signed [31:0] shifted_state_out108_0 = reservoir_state[108] <<< 0;
wire signed [31:0] shifted_state_out108_3 = reservoir_state[108] <<< 3;
wire signed [31:0] shifted_state_out109_2 = reservoir_state[109] <<< 2;
wire signed [31:0] shifted_state_out109_3 = reservoir_state[109] <<< 3;
wire signed [31:0] shifted_state_out109_4 = reservoir_state[109] <<< 4;
wire signed [31:0] shifted_state_out109_5 = reservoir_state[109] <<< 5;
wire signed [31:0] shifted_state_out109_6 = reservoir_state[109] <<< 6;
wire signed [31:0] shifted_state_out109_7 = reservoir_state[109] <<< 7;
wire signed [31:0] shifted_state_out111_0 = reservoir_state[111] <<< 0;
wire signed [31:0] shifted_state_out111_1 = reservoir_state[111] <<< 1;
wire signed [31:0] shifted_state_out112_1 = reservoir_state[112] <<< 1;
wire signed [31:0] shifted_state_out112_3 = reservoir_state[112] <<< 3;
wire signed [31:0] shifted_state_out112_4 = reservoir_state[112] <<< 4;
wire signed [31:0] shifted_state_out112_5 = reservoir_state[112] <<< 5;
wire signed [31:0] shifted_state_out112_6 = reservoir_state[112] <<< 6;
wire signed [31:0] shifted_state_out112_7 = reservoir_state[112] <<< 7;
wire signed [31:0] shifted_state_out113_1 = reservoir_state[113] <<< 1;
wire signed [31:0] shifted_state_out113_3 = reservoir_state[113] <<< 3;
wire signed [31:0] shifted_state_out113_4 = reservoir_state[113] <<< 4;
wire signed [31:0] shifted_state_out113_5 = reservoir_state[113] <<< 5;
wire signed [31:0] shifted_state_out113_6 = reservoir_state[113] <<< 6;
wire signed [31:0] shifted_state_out113_7 = reservoir_state[113] <<< 7;
wire signed [31:0] shifted_state_out114_0 = reservoir_state[114] <<< 0;
wire signed [31:0] shifted_state_out114_2 = reservoir_state[114] <<< 2;
wire signed [31:0] shifted_state_out114_3 = reservoir_state[114] <<< 3;
wire signed [31:0] shifted_state_out114_4 = reservoir_state[114] <<< 4;
wire signed [31:0] shifted_state_out114_5 = reservoir_state[114] <<< 5;
wire signed [31:0] shifted_state_out114_6 = reservoir_state[114] <<< 6;
wire signed [31:0] shifted_state_out114_7 = reservoir_state[114] <<< 7;
wire signed [31:0] shifted_state_out115_1 = reservoir_state[115] <<< 1;
wire signed [31:0] shifted_state_out115_3 = reservoir_state[115] <<< 3;
wire signed [31:0] shifted_state_out115_4 = reservoir_state[115] <<< 4;
wire signed [31:0] shifted_state_out115_5 = reservoir_state[115] <<< 5;
wire signed [31:0] shifted_state_out115_6 = reservoir_state[115] <<< 6;
wire signed [31:0] shifted_state_out115_7 = reservoir_state[115] <<< 7;
wire signed [31:0] shifted_state_out116_0 = reservoir_state[116] <<< 0;
wire signed [31:0] shifted_state_out117_0 = reservoir_state[117] <<< 0;
wire signed [31:0] shifted_state_out117_2 = reservoir_state[117] <<< 2;
wire signed [31:0] shifted_state_out118_1 = reservoir_state[118] <<< 1;
wire signed [31:0] shifted_state_out118_2 = reservoir_state[118] <<< 2;
wire signed [31:0] shifted_state_out119_0 = reservoir_state[119] <<< 0;
wire signed [31:0] shifted_state_out119_1 = reservoir_state[119] <<< 1;
wire signed [31:0] shifted_state_out119_2 = reservoir_state[119] <<< 2;
wire signed [31:0] shifted_state_out119_3 = reservoir_state[119] <<< 3;
wire signed [31:0] shifted_state_out119_4 = reservoir_state[119] <<< 4;
wire signed [31:0] shifted_state_out119_5 = reservoir_state[119] <<< 5;
wire signed [31:0] shifted_state_out119_6 = reservoir_state[119] <<< 6;
wire signed [31:0] shifted_state_out119_7 = reservoir_state[119] <<< 7;
wire signed [31:0] shifted_state_out120_0 = reservoir_state[120] <<< 0;
wire signed [31:0] shifted_state_out120_1 = reservoir_state[120] <<< 1;
wire signed [31:0] shifted_state_out120_3 = reservoir_state[120] <<< 3;
wire signed [31:0] shifted_state_out120_4 = reservoir_state[120] <<< 4;
wire signed [31:0] shifted_state_out120_5 = reservoir_state[120] <<< 5;
wire signed [31:0] shifted_state_out120_6 = reservoir_state[120] <<< 6;
wire signed [31:0] shifted_state_out120_7 = reservoir_state[120] <<< 7;
wire signed [31:0] shifted_state_out121_0 = reservoir_state[121] <<< 0;
wire signed [31:0] shifted_state_out121_2 = reservoir_state[121] <<< 2;
wire signed [31:0] shifted_state_out121_3 = reservoir_state[121] <<< 3;
wire signed [31:0] shifted_state_out121_4 = reservoir_state[121] <<< 4;
wire signed [31:0] shifted_state_out121_5 = reservoir_state[121] <<< 5;
wire signed [31:0] shifted_state_out121_6 = reservoir_state[121] <<< 6;
wire signed [31:0] shifted_state_out121_7 = reservoir_state[121] <<< 7;
wire signed [31:0] shifted_state_out122_0 = reservoir_state[122] <<< 0;
wire signed [31:0] shifted_state_out122_2 = reservoir_state[122] <<< 2;
wire signed [31:0] shifted_state_out123_0 = reservoir_state[123] <<< 0;
wire signed [31:0] shifted_state_out123_1 = reservoir_state[123] <<< 1;
wire signed [31:0] shifted_state_out124_1 = reservoir_state[124] <<< 1;
wire signed [31:0] shifted_state_out124_2 = reservoir_state[124] <<< 2;
wire signed [31:0] shifted_state_out124_3 = reservoir_state[124] <<< 3;
wire signed [31:0] shifted_state_out124_4 = reservoir_state[124] <<< 4;
wire signed [31:0] shifted_state_out124_5 = reservoir_state[124] <<< 5;
wire signed [31:0] shifted_state_out124_6 = reservoir_state[124] <<< 6;
wire signed [31:0] shifted_state_out124_7 = reservoir_state[124] <<< 7;
wire signed [31:0] shifted_state_out125_0 = reservoir_state[125] <<< 0;
wire signed [31:0] shifted_state_out125_1 = reservoir_state[125] <<< 1;
wire signed [31:0] shifted_state_out125_2 = reservoir_state[125] <<< 2;
wire signed [31:0] shifted_state_out125_3 = reservoir_state[125] <<< 3;
wire signed [31:0] shifted_state_out125_4 = reservoir_state[125] <<< 4;
wire signed [31:0] shifted_state_out125_5 = reservoir_state[125] <<< 5;
wire signed [31:0] shifted_state_out125_6 = reservoir_state[125] <<< 6;
wire signed [31:0] shifted_state_out125_7 = reservoir_state[125] <<< 7;
wire signed [31:0] shifted_state_out126_1 = reservoir_state[126] <<< 1;
wire signed [31:0] shifted_state_out126_2 = reservoir_state[126] <<< 2;
wire signed [31:0] shifted_state_out127_1 = reservoir_state[127] <<< 1;
wire signed [31:0] shifted_state_out128_0 = reservoir_state[128] <<< 0;
wire signed [31:0] shifted_state_out128_1 = reservoir_state[128] <<< 1;
wire signed [31:0] shifted_state_out129_1 = reservoir_state[129] <<< 1;
wire signed [31:0] shifted_state_out129_2 = reservoir_state[129] <<< 2;
wire signed [31:0] shifted_state_out129_3 = reservoir_state[129] <<< 3;
wire signed [31:0] shifted_state_out129_4 = reservoir_state[129] <<< 4;
wire signed [31:0] shifted_state_out129_5 = reservoir_state[129] <<< 5;
wire signed [31:0] shifted_state_out129_6 = reservoir_state[129] <<< 6;
wire signed [31:0] shifted_state_out129_7 = reservoir_state[129] <<< 7;
wire signed [31:0] shifted_state_out131_0 = reservoir_state[131] <<< 0;
wire signed [31:0] shifted_state_out132_0 = reservoir_state[132] <<< 0;
wire signed [31:0] shifted_state_out133_0 = reservoir_state[133] <<< 0;
wire signed [31:0] shifted_state_out133_1 = reservoir_state[133] <<< 1;
wire signed [31:0] shifted_state_out134_1 = reservoir_state[134] <<< 1;
wire signed [31:0] shifted_state_out134_2 = reservoir_state[134] <<< 2;
wire signed [31:0] shifted_state_out135_0 = reservoir_state[135] <<< 0;
wire signed [31:0] shifted_state_out135_1 = reservoir_state[135] <<< 1;
wire signed [31:0] shifted_state_out135_2 = reservoir_state[135] <<< 2;
wire signed [31:0] shifted_state_out135_3 = reservoir_state[135] <<< 3;
wire signed [31:0] shifted_state_out135_4 = reservoir_state[135] <<< 4;
wire signed [31:0] shifted_state_out135_5 = reservoir_state[135] <<< 5;
wire signed [31:0] shifted_state_out135_6 = reservoir_state[135] <<< 6;
wire signed [31:0] shifted_state_out135_7 = reservoir_state[135] <<< 7;
wire signed [31:0] shifted_state_out137_0 = reservoir_state[137] <<< 0;
wire signed [31:0] shifted_state_out137_2 = reservoir_state[137] <<< 2;
wire signed [31:0] shifted_state_out138_2 = reservoir_state[138] <<< 2;
wire signed [31:0] shifted_state_out138_3 = reservoir_state[138] <<< 3;
wire signed [31:0] shifted_state_out138_4 = reservoir_state[138] <<< 4;
wire signed [31:0] shifted_state_out138_5 = reservoir_state[138] <<< 5;
wire signed [31:0] shifted_state_out138_6 = reservoir_state[138] <<< 6;
wire signed [31:0] shifted_state_out138_7 = reservoir_state[138] <<< 7;
wire signed [31:0] shifted_state_out139_0 = reservoir_state[139] <<< 0;
wire signed [31:0] shifted_state_out139_1 = reservoir_state[139] <<< 1;
wire signed [31:0] shifted_state_out139_2 = reservoir_state[139] <<< 2;
wire signed [31:0] shifted_state_out139_3 = reservoir_state[139] <<< 3;
wire signed [31:0] shifted_state_out139_4 = reservoir_state[139] <<< 4;
wire signed [31:0] shifted_state_out139_5 = reservoir_state[139] <<< 5;
wire signed [31:0] shifted_state_out139_6 = reservoir_state[139] <<< 6;
wire signed [31:0] shifted_state_out139_7 = reservoir_state[139] <<< 7;
wire signed [31:0] shifted_state_out140_0 = reservoir_state[140] <<< 0;
wire signed [31:0] shifted_state_out140_1 = reservoir_state[140] <<< 1;
wire signed [31:0] shifted_state_out140_2 = reservoir_state[140] <<< 2;
wire signed [31:0] shifted_state_out140_3 = reservoir_state[140] <<< 3;
wire signed [31:0] shifted_state_out140_4 = reservoir_state[140] <<< 4;
wire signed [31:0] shifted_state_out140_5 = reservoir_state[140] <<< 5;
wire signed [31:0] shifted_state_out140_6 = reservoir_state[140] <<< 6;
wire signed [31:0] shifted_state_out140_7 = reservoir_state[140] <<< 7;
wire signed [31:0] shifted_state_out141_2 = reservoir_state[141] <<< 2;
wire signed [31:0] shifted_state_out142_1 = reservoir_state[142] <<< 1;
wire signed [31:0] shifted_state_out142_2 = reservoir_state[142] <<< 2;
wire signed [31:0] shifted_state_out142_3 = reservoir_state[142] <<< 3;
wire signed [31:0] shifted_state_out142_4 = reservoir_state[142] <<< 4;
wire signed [31:0] shifted_state_out142_5 = reservoir_state[142] <<< 5;
wire signed [31:0] shifted_state_out142_6 = reservoir_state[142] <<< 6;
wire signed [31:0] shifted_state_out142_7 = reservoir_state[142] <<< 7;
wire signed [31:0] shifted_state_out143_0 = reservoir_state[143] <<< 0;
wire signed [31:0] shifted_state_out143_1 = reservoir_state[143] <<< 1;
wire signed [31:0] shifted_state_out143_2 = reservoir_state[143] <<< 2;
wire signed [31:0] shifted_state_out143_3 = reservoir_state[143] <<< 3;
wire signed [31:0] shifted_state_out143_4 = reservoir_state[143] <<< 4;
wire signed [31:0] shifted_state_out143_5 = reservoir_state[143] <<< 5;
wire signed [31:0] shifted_state_out143_6 = reservoir_state[143] <<< 6;
wire signed [31:0] shifted_state_out143_7 = reservoir_state[143] <<< 7;
wire signed [31:0] shifted_state_out144_2 = reservoir_state[144] <<< 2;
wire signed [31:0] shifted_state_out144_3 = reservoir_state[144] <<< 3;
wire signed [31:0] shifted_state_out144_4 = reservoir_state[144] <<< 4;
wire signed [31:0] shifted_state_out144_5 = reservoir_state[144] <<< 5;
wire signed [31:0] shifted_state_out144_6 = reservoir_state[144] <<< 6;
wire signed [31:0] shifted_state_out144_7 = reservoir_state[144] <<< 7;
wire signed [31:0] shifted_state_out145_0 = reservoir_state[145] <<< 0;
wire signed [31:0] shifted_state_out145_1 = reservoir_state[145] <<< 1;
wire signed [31:0] shifted_state_out145_2 = reservoir_state[145] <<< 2;
wire signed [31:0] shifted_state_out145_3 = reservoir_state[145] <<< 3;
wire signed [31:0] shifted_state_out145_4 = reservoir_state[145] <<< 4;
wire signed [31:0] shifted_state_out145_5 = reservoir_state[145] <<< 5;
wire signed [31:0] shifted_state_out145_6 = reservoir_state[145] <<< 6;
wire signed [31:0] shifted_state_out145_7 = reservoir_state[145] <<< 7;
wire signed [31:0] shifted_state_out146_0 = reservoir_state[146] <<< 0;
wire signed [31:0] shifted_state_out146_1 = reservoir_state[146] <<< 1;
wire signed [31:0] shifted_state_out146_3 = reservoir_state[146] <<< 3;
wire signed [31:0] shifted_state_out146_4 = reservoir_state[146] <<< 4;
wire signed [31:0] shifted_state_out146_5 = reservoir_state[146] <<< 5;
wire signed [31:0] shifted_state_out146_6 = reservoir_state[146] <<< 6;
wire signed [31:0] shifted_state_out146_7 = reservoir_state[146] <<< 7;
wire signed [31:0] shifted_state_out147_0 = reservoir_state[147] <<< 0;
wire signed [31:0] shifted_state_out147_1 = reservoir_state[147] <<< 1;
wire signed [31:0] shifted_state_out147_2 = reservoir_state[147] <<< 2;
wire signed [31:0] shifted_state_out148_1 = reservoir_state[148] <<< 1;
wire signed [31:0] shifted_state_out149_1 = reservoir_state[149] <<< 1;
wire signed [31:0] shifted_state_out149_3 = reservoir_state[149] <<< 3;
wire signed [31:0] shifted_state_out150_0 = reservoir_state[150] <<< 0;
wire signed [31:0] shifted_state_out150_2 = reservoir_state[150] <<< 2;
wire signed [31:0] shifted_state_out150_3 = reservoir_state[150] <<< 3;
wire signed [31:0] shifted_state_out150_4 = reservoir_state[150] <<< 4;
wire signed [31:0] shifted_state_out150_5 = reservoir_state[150] <<< 5;
wire signed [31:0] shifted_state_out150_6 = reservoir_state[150] <<< 6;
wire signed [31:0] shifted_state_out150_7 = reservoir_state[150] <<< 7;
wire signed [31:0] shifted_state_out151_1 = reservoir_state[151] <<< 1;
wire signed [31:0] shifted_state_out151_2 = reservoir_state[151] <<< 2;
wire signed [31:0] shifted_state_out151_3 = reservoir_state[151] <<< 3;
wire signed [31:0] shifted_state_out151_4 = reservoir_state[151] <<< 4;
wire signed [31:0] shifted_state_out151_5 = reservoir_state[151] <<< 5;
wire signed [31:0] shifted_state_out151_6 = reservoir_state[151] <<< 6;
wire signed [31:0] shifted_state_out151_7 = reservoir_state[151] <<< 7;
wire signed [31:0] shifted_state_out152_1 = reservoir_state[152] <<< 1;
wire signed [31:0] shifted_state_out152_2 = reservoir_state[152] <<< 2;
wire signed [31:0] shifted_state_out152_3 = reservoir_state[152] <<< 3;
wire signed [31:0] shifted_state_out152_4 = reservoir_state[152] <<< 4;
wire signed [31:0] shifted_state_out152_5 = reservoir_state[152] <<< 5;
wire signed [31:0] shifted_state_out152_6 = reservoir_state[152] <<< 6;
wire signed [31:0] shifted_state_out152_7 = reservoir_state[152] <<< 7;
wire signed [31:0] shifted_state_out153_0 = reservoir_state[153] <<< 0;
wire signed [31:0] shifted_state_out153_2 = reservoir_state[153] <<< 2;
wire signed [31:0] shifted_state_out153_3 = reservoir_state[153] <<< 3;
wire signed [31:0] shifted_state_out153_4 = reservoir_state[153] <<< 4;
wire signed [31:0] shifted_state_out153_5 = reservoir_state[153] <<< 5;
wire signed [31:0] shifted_state_out153_6 = reservoir_state[153] <<< 6;
wire signed [31:0] shifted_state_out153_7 = reservoir_state[153] <<< 7;
wire signed [31:0] shifted_state_out154_1 = reservoir_state[154] <<< 1;
wire signed [31:0] shifted_state_out154_2 = reservoir_state[154] <<< 2;
wire signed [31:0] shifted_state_out154_3 = reservoir_state[154] <<< 3;
wire signed [31:0] shifted_state_out154_4 = reservoir_state[154] <<< 4;
wire signed [31:0] shifted_state_out154_5 = reservoir_state[154] <<< 5;
wire signed [31:0] shifted_state_out154_6 = reservoir_state[154] <<< 6;
wire signed [31:0] shifted_state_out154_7 = reservoir_state[154] <<< 7;
wire signed [31:0] shifted_state_out155_0 = reservoir_state[155] <<< 0;
wire signed [31:0] shifted_state_out155_7 = reservoir_state[155] <<< 7;
wire signed [31:0] shifted_state_out156_3 = reservoir_state[156] <<< 3;
wire signed [31:0] shifted_state_out156_4 = reservoir_state[156] <<< 4;
wire signed [31:0] shifted_state_out156_5 = reservoir_state[156] <<< 5;
wire signed [31:0] shifted_state_out156_6 = reservoir_state[156] <<< 6;
wire signed [31:0] shifted_state_out156_7 = reservoir_state[156] <<< 7;
wire signed [31:0] shifted_state_out157_1 = reservoir_state[157] <<< 1;
wire signed [31:0] shifted_state_out157_2 = reservoir_state[157] <<< 2;
wire signed [31:0] shifted_state_out157_3 = reservoir_state[157] <<< 3;
wire signed [31:0] shifted_state_out157_4 = reservoir_state[157] <<< 4;
wire signed [31:0] shifted_state_out157_5 = reservoir_state[157] <<< 5;
wire signed [31:0] shifted_state_out157_6 = reservoir_state[157] <<< 6;
wire signed [31:0] shifted_state_out157_7 = reservoir_state[157] <<< 7;
wire signed [31:0] shifted_state_out158_2 = reservoir_state[158] <<< 2;
wire signed [31:0] shifted_state_out158_3 = reservoir_state[158] <<< 3;
wire signed [31:0] shifted_state_out158_4 = reservoir_state[158] <<< 4;
wire signed [31:0] shifted_state_out158_5 = reservoir_state[158] <<< 5;
wire signed [31:0] shifted_state_out158_6 = reservoir_state[158] <<< 6;
wire signed [31:0] shifted_state_out158_7 = reservoir_state[158] <<< 7;
wire signed [31:0] shifted_state_out159_0 = reservoir_state[159] <<< 0;
wire signed [31:0] shifted_state_out159_2 = reservoir_state[159] <<< 2;
wire signed [31:0] shifted_state_out160_2 = reservoir_state[160] <<< 2;
wire signed [31:0] shifted_state_out160_3 = reservoir_state[160] <<< 3;
wire signed [31:0] shifted_state_out160_4 = reservoir_state[160] <<< 4;
wire signed [31:0] shifted_state_out160_5 = reservoir_state[160] <<< 5;
wire signed [31:0] shifted_state_out160_6 = reservoir_state[160] <<< 6;
wire signed [31:0] shifted_state_out160_7 = reservoir_state[160] <<< 7;
wire signed [31:0] shifted_state_out161_0 = reservoir_state[161] <<< 0;
wire signed [31:0] shifted_state_out161_1 = reservoir_state[161] <<< 1;
wire signed [31:0] shifted_state_out161_2 = reservoir_state[161] <<< 2;
wire signed [31:0] shifted_state_out161_3 = reservoir_state[161] <<< 3;
wire signed [31:0] shifted_state_out161_4 = reservoir_state[161] <<< 4;
wire signed [31:0] shifted_state_out161_5 = reservoir_state[161] <<< 5;
wire signed [31:0] shifted_state_out161_6 = reservoir_state[161] <<< 6;
wire signed [31:0] shifted_state_out161_7 = reservoir_state[161] <<< 7;
wire signed [31:0] shifted_state_out162_1 = reservoir_state[162] <<< 1;
wire signed [31:0] shifted_state_out162_2 = reservoir_state[162] <<< 2;
wire signed [31:0] shifted_state_out162_3 = reservoir_state[162] <<< 3;
wire signed [31:0] shifted_state_out162_4 = reservoir_state[162] <<< 4;
wire signed [31:0] shifted_state_out162_5 = reservoir_state[162] <<< 5;
wire signed [31:0] shifted_state_out162_6 = reservoir_state[162] <<< 6;
wire signed [31:0] shifted_state_out162_7 = reservoir_state[162] <<< 7;
wire signed [31:0] shifted_state_out164_0 = reservoir_state[164] <<< 0;
wire signed [31:0] shifted_state_out164_3 = reservoir_state[164] <<< 3;
wire signed [31:0] shifted_state_out164_4 = reservoir_state[164] <<< 4;
wire signed [31:0] shifted_state_out164_5 = reservoir_state[164] <<< 5;
wire signed [31:0] shifted_state_out164_6 = reservoir_state[164] <<< 6;
wire signed [31:0] shifted_state_out164_7 = reservoir_state[164] <<< 7;
wire signed [31:0] shifted_state_out165_0 = reservoir_state[165] <<< 0;
wire signed [31:0] shifted_state_out165_2 = reservoir_state[165] <<< 2;
wire signed [31:0] shifted_state_out166_0 = reservoir_state[166] <<< 0;
wire signed [31:0] shifted_state_out166_1 = reservoir_state[166] <<< 1;
wire signed [31:0] shifted_state_out166_3 = reservoir_state[166] <<< 3;
wire signed [31:0] shifted_state_out166_4 = reservoir_state[166] <<< 4;
wire signed [31:0] shifted_state_out166_5 = reservoir_state[166] <<< 5;
wire signed [31:0] shifted_state_out166_6 = reservoir_state[166] <<< 6;
wire signed [31:0] shifted_state_out166_7 = reservoir_state[166] <<< 7;
wire signed [31:0] shifted_state_out167_1 = reservoir_state[167] <<< 1;
wire signed [31:0] shifted_state_out167_2 = reservoir_state[167] <<< 2;
wire signed [31:0] shifted_state_out167_3 = reservoir_state[167] <<< 3;
wire signed [31:0] shifted_state_out167_4 = reservoir_state[167] <<< 4;
wire signed [31:0] shifted_state_out167_5 = reservoir_state[167] <<< 5;
wire signed [31:0] shifted_state_out167_6 = reservoir_state[167] <<< 6;
wire signed [31:0] shifted_state_out167_7 = reservoir_state[167] <<< 7;
wire signed [31:0] shifted_state_out169_1 = reservoir_state[169] <<< 1;
wire signed [31:0] shifted_state_out170_0 = reservoir_state[170] <<< 0;
wire signed [31:0] shifted_state_out170_2 = reservoir_state[170] <<< 2;
wire signed [31:0] shifted_state_out171_2 = reservoir_state[171] <<< 2;
wire signed [31:0] shifted_state_out172_1 = reservoir_state[172] <<< 1;
wire signed [31:0] shifted_state_out173_1 = reservoir_state[173] <<< 1;
wire signed [31:0] shifted_state_out173_2 = reservoir_state[173] <<< 2;
wire signed [31:0] shifted_state_out174_3 = reservoir_state[174] <<< 3;
wire signed [31:0] shifted_state_out174_4 = reservoir_state[174] <<< 4;
wire signed [31:0] shifted_state_out174_5 = reservoir_state[174] <<< 5;
wire signed [31:0] shifted_state_out174_6 = reservoir_state[174] <<< 6;
wire signed [31:0] shifted_state_out174_7 = reservoir_state[174] <<< 7;
wire signed [31:0] shifted_state_out175_0 = reservoir_state[175] <<< 0;
wire signed [31:0] shifted_state_out175_1 = reservoir_state[175] <<< 1;
wire signed [31:0] shifted_state_out176_0 = reservoir_state[176] <<< 0;
wire signed [31:0] shifted_state_out176_1 = reservoir_state[176] <<< 1;
wire signed [31:0] shifted_state_out177_1 = reservoir_state[177] <<< 1;
wire signed [31:0] shifted_state_out177_2 = reservoir_state[177] <<< 2;
wire signed [31:0] shifted_state_out178_0 = reservoir_state[178] <<< 0;
wire signed [31:0] shifted_state_out178_2 = reservoir_state[178] <<< 2;
wire signed [31:0] shifted_state_out178_4 = reservoir_state[178] <<< 4;
wire signed [31:0] shifted_state_out178_5 = reservoir_state[178] <<< 5;
wire signed [31:0] shifted_state_out178_6 = reservoir_state[178] <<< 6;
wire signed [31:0] shifted_state_out178_7 = reservoir_state[178] <<< 7;
wire signed [31:0] shifted_state_out179_3 = reservoir_state[179] <<< 3;
wire signed [31:0] shifted_state_out179_4 = reservoir_state[179] <<< 4;
wire signed [31:0] shifted_state_out179_5 = reservoir_state[179] <<< 5;
wire signed [31:0] shifted_state_out179_6 = reservoir_state[179] <<< 6;
wire signed [31:0] shifted_state_out179_7 = reservoir_state[179] <<< 7;
wire signed [31:0] shifted_state_out180_0 = reservoir_state[180] <<< 0;
wire signed [31:0] shifted_state_out180_1 = reservoir_state[180] <<< 1;
wire signed [31:0] shifted_state_out181_3 = reservoir_state[181] <<< 3;
wire signed [31:0] shifted_state_out181_4 = reservoir_state[181] <<< 4;
wire signed [31:0] shifted_state_out181_5 = reservoir_state[181] <<< 5;
wire signed [31:0] shifted_state_out181_6 = reservoir_state[181] <<< 6;
wire signed [31:0] shifted_state_out181_7 = reservoir_state[181] <<< 7;
wire signed [31:0] shifted_state_out182_0 = reservoir_state[182] <<< 0;
wire signed [31:0] shifted_state_out182_3 = reservoir_state[182] <<< 3;
wire signed [31:0] shifted_state_out183_0 = reservoir_state[183] <<< 0;
wire signed [31:0] shifted_state_out183_2 = reservoir_state[183] <<< 2;
wire signed [31:0] shifted_state_out183_3 = reservoir_state[183] <<< 3;
wire signed [31:0] shifted_state_out183_4 = reservoir_state[183] <<< 4;
wire signed [31:0] shifted_state_out183_5 = reservoir_state[183] <<< 5;
wire signed [31:0] shifted_state_out183_6 = reservoir_state[183] <<< 6;
wire signed [31:0] shifted_state_out183_7 = reservoir_state[183] <<< 7;
wire signed [31:0] shifted_state_out184_0 = reservoir_state[184] <<< 0;
wire signed [31:0] shifted_state_out184_1 = reservoir_state[184] <<< 1;
wire signed [31:0] shifted_state_out185_0 = reservoir_state[185] <<< 0;
wire signed [31:0] shifted_state_out185_1 = reservoir_state[185] <<< 1;
wire signed [31:0] shifted_state_out185_2 = reservoir_state[185] <<< 2;
wire signed [31:0] shifted_state_out186_2 = reservoir_state[186] <<< 2;
wire signed [31:0] shifted_state_out186_3 = reservoir_state[186] <<< 3;
wire signed [31:0] shifted_state_out186_4 = reservoir_state[186] <<< 4;
wire signed [31:0] shifted_state_out186_5 = reservoir_state[186] <<< 5;
wire signed [31:0] shifted_state_out186_6 = reservoir_state[186] <<< 6;
wire signed [31:0] shifted_state_out186_7 = reservoir_state[186] <<< 7;
wire signed [31:0] shifted_state_out187_1 = reservoir_state[187] <<< 1;
wire signed [31:0] shifted_state_out188_0 = reservoir_state[188] <<< 0;
wire signed [31:0] shifted_state_out188_2 = reservoir_state[188] <<< 2;
wire signed [31:0] shifted_state_out188_3 = reservoir_state[188] <<< 3;
wire signed [31:0] shifted_state_out188_4 = reservoir_state[188] <<< 4;
wire signed [31:0] shifted_state_out188_5 = reservoir_state[188] <<< 5;
wire signed [31:0] shifted_state_out188_6 = reservoir_state[188] <<< 6;
wire signed [31:0] shifted_state_out188_7 = reservoir_state[188] <<< 7;
wire signed [31:0] shifted_state_out189_1 = reservoir_state[189] <<< 1;
wire signed [31:0] shifted_state_out190_1 = reservoir_state[190] <<< 1;
wire signed [31:0] shifted_state_out190_2 = reservoir_state[190] <<< 2;
wire signed [31:0] shifted_state_out190_3 = reservoir_state[190] <<< 3;
wire signed [31:0] shifted_state_out190_4 = reservoir_state[190] <<< 4;
wire signed [31:0] shifted_state_out190_5 = reservoir_state[190] <<< 5;
wire signed [31:0] shifted_state_out190_6 = reservoir_state[190] <<< 6;
wire signed [31:0] shifted_state_out190_7 = reservoir_state[190] <<< 7;
wire signed [31:0] shifted_state_out191_1 = reservoir_state[191] <<< 1;
wire signed [31:0] shifted_state_out192_0 = reservoir_state[192] <<< 0;
wire signed [31:0] shifted_state_out193_0 = reservoir_state[193] <<< 0;
wire signed [31:0] shifted_state_out193_2 = reservoir_state[193] <<< 2;
wire signed [31:0] shifted_state_out193_3 = reservoir_state[193] <<< 3;
wire signed [31:0] shifted_state_out193_4 = reservoir_state[193] <<< 4;
wire signed [31:0] shifted_state_out193_5 = reservoir_state[193] <<< 5;
wire signed [31:0] shifted_state_out193_6 = reservoir_state[193] <<< 6;
wire signed [31:0] shifted_state_out193_7 = reservoir_state[193] <<< 7;
wire signed [31:0] shifted_state_out194_0 = reservoir_state[194] <<< 0;
wire signed [31:0] shifted_state_out194_1 = reservoir_state[194] <<< 1;
wire signed [31:0] shifted_state_out194_2 = reservoir_state[194] <<< 2;
wire signed [31:0] shifted_state_out194_3 = reservoir_state[194] <<< 3;
wire signed [31:0] shifted_state_out194_4 = reservoir_state[194] <<< 4;
wire signed [31:0] shifted_state_out194_5 = reservoir_state[194] <<< 5;
wire signed [31:0] shifted_state_out194_6 = reservoir_state[194] <<< 6;
wire signed [31:0] shifted_state_out194_7 = reservoir_state[194] <<< 7;
wire signed [31:0] shifted_state_out195_0 = reservoir_state[195] <<< 0;
wire signed [31:0] shifted_state_out195_1 = reservoir_state[195] <<< 1;
wire signed [31:0] shifted_state_out195_2 = reservoir_state[195] <<< 2;
wire signed [31:0] shifted_state_out195_3 = reservoir_state[195] <<< 3;
wire signed [31:0] shifted_state_out195_4 = reservoir_state[195] <<< 4;
wire signed [31:0] shifted_state_out195_5 = reservoir_state[195] <<< 5;
wire signed [31:0] shifted_state_out195_6 = reservoir_state[195] <<< 6;
wire signed [31:0] shifted_state_out195_7 = reservoir_state[195] <<< 7;
wire signed [31:0] shifted_state_out196_1 = reservoir_state[196] <<< 1;
wire signed [31:0] shifted_state_out196_2 = reservoir_state[196] <<< 2;
wire signed [31:0] shifted_state_out196_3 = reservoir_state[196] <<< 3;
wire signed [31:0] shifted_state_out196_4 = reservoir_state[196] <<< 4;
wire signed [31:0] shifted_state_out196_5 = reservoir_state[196] <<< 5;
wire signed [31:0] shifted_state_out196_6 = reservoir_state[196] <<< 6;
wire signed [31:0] shifted_state_out196_7 = reservoir_state[196] <<< 7;
wire signed [31:0] shifted_state_out197_1 = reservoir_state[197] <<< 1;
wire signed [31:0] shifted_state_out197_2 = reservoir_state[197] <<< 2;
wire signed [31:0] shifted_state_out197_3 = reservoir_state[197] <<< 3;
wire signed [31:0] shifted_state_out197_4 = reservoir_state[197] <<< 4;
wire signed [31:0] shifted_state_out197_5 = reservoir_state[197] <<< 5;
wire signed [31:0] shifted_state_out197_6 = reservoir_state[197] <<< 6;
wire signed [31:0] shifted_state_out197_7 = reservoir_state[197] <<< 7;
wire signed [31:0] shifted_state_out198_0 = reservoir_state[198] <<< 0;
wire signed [31:0] shifted_state_out198_1 = reservoir_state[198] <<< 1;
wire signed [31:0] shifted_state_out198_3 = reservoir_state[198] <<< 3;
wire signed [31:0] shifted_state_out198_4 = reservoir_state[198] <<< 4;
wire signed [31:0] shifted_state_out198_5 = reservoir_state[198] <<< 5;
wire signed [31:0] shifted_state_out198_6 = reservoir_state[198] <<< 6;
wire signed [31:0] shifted_state_out198_7 = reservoir_state[198] <<< 7;
wire signed [31:0] shifted_state_out199_0 = reservoir_state[199] <<< 0;
wire signed [31:0] shifted_state_out199_1 = reservoir_state[199] <<< 1;
wire signed [31:0] shifted_state_out199_3 = reservoir_state[199] <<< 3;
wire signed [31:0] shifted_state_out199_4 = reservoir_state[199] <<< 4;
wire signed [31:0] shifted_state_out199_5 = reservoir_state[199] <<< 5;
wire signed [31:0] shifted_state_out199_6 = reservoir_state[199] <<< 6;
wire signed [31:0] shifted_state_out199_7 = reservoir_state[199] <<< 7;
wire signed [31:0] shifted_input0 = input_data <<< 0;
wire signed [31:0] shifted_input1 = input_data <<< 1;
wire signed [31:0] shifted_input2 = input_data <<< 2;
wire signed [31:0] shifted_input3 = input_data <<< 3;
wire signed [31:0] shifted_input4 = input_data <<< 4;
wire signed [31:0] shifted_input5 = input_data <<< 5;
wire signed [31:0] shifted_input6 = input_data <<< 6;
wire signed [31:0] shifted_input7 = input_data <<< 7;

  // ESN logic
  always @(posedge clk) begin

      input_sum_parallel[0] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[1] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[2] = 0;
      input_sum_parallel[3] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[4] = shifted_input7;
      input_sum_parallel[5] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[6] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[7] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[8] = shifted_input7;
      input_sum_parallel[9] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[10] = shifted_input7;
      input_sum_parallel[11] = 0;
      input_sum_parallel[12] = shifted_input7;
      input_sum_parallel[13] = shifted_input7;
      input_sum_parallel[14] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[15] = 0;
      input_sum_parallel[16] = shifted_input7;
      input_sum_parallel[17] = shifted_input7;
      input_sum_parallel[18] = shifted_input7;
      input_sum_parallel[19] = shifted_input7;
      input_sum_parallel[20] = 0;
      input_sum_parallel[21] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[22] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[23] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[24] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[25] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[26] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[27] = shifted_input7;
      input_sum_parallel[28] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[29] = shifted_input7;
      input_sum_parallel[30] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[31] = shifted_input7;
      input_sum_parallel[32] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[33] = 0;
      input_sum_parallel[34] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[35] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[36] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[37] = shifted_input7;
      input_sum_parallel[38] = shifted_input7;
      input_sum_parallel[39] = shifted_input7;
      input_sum_parallel[40] = 0;
      input_sum_parallel[41] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[42] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[43] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[44] = shifted_input7;
      input_sum_parallel[45] = shifted_input7;
      input_sum_parallel[46] = shifted_input7;
      input_sum_parallel[47] = shifted_input7;
      input_sum_parallel[48] = 0;
      input_sum_parallel[49] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[50] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[51] = shifted_input7;
      input_sum_parallel[52] = shifted_input7;
      input_sum_parallel[53] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[54] = shifted_input7;
      input_sum_parallel[55] = shifted_input7;
      input_sum_parallel[56] = shifted_input7;
      input_sum_parallel[57] = shifted_input7;
      input_sum_parallel[58] = shifted_input7;
      input_sum_parallel[59] = 0;
      input_sum_parallel[60] = shifted_input7;
      input_sum_parallel[61] = shifted_input7;
      input_sum_parallel[62] = shifted_input7;
      input_sum_parallel[63] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[64] = shifted_input7;
      input_sum_parallel[65] = shifted_input7;
      input_sum_parallel[66] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[67] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[68] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[69] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[70] = shifted_input7;
      input_sum_parallel[71] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[72] = shifted_input7;
      input_sum_parallel[73] = shifted_input7;
      input_sum_parallel[74] = shifted_input7;
      input_sum_parallel[75] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[76] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[77] = shifted_input7;
      input_sum_parallel[78] = shifted_input7;
      input_sum_parallel[79] = shifted_input7;
      input_sum_parallel[80] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[81] = shifted_input7;
      input_sum_parallel[82] = shifted_input7;
      input_sum_parallel[83] = shifted_input7;
      input_sum_parallel[84] = shifted_input7;
      input_sum_parallel[85] = shifted_input7;
      input_sum_parallel[86] = 0;
      input_sum_parallel[87] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[88] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[89] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[90] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[91] = shifted_input7;
      input_sum_parallel[92] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[93] = shifted_input7;
      input_sum_parallel[94] = shifted_input7;
      input_sum_parallel[95] = 0;
      input_sum_parallel[96] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[97] = shifted_input7;
      input_sum_parallel[98] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[99] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[100] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[101] = 0;
      input_sum_parallel[102] = shifted_input7;
      input_sum_parallel[103] = 0;
      input_sum_parallel[104] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[105] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[106] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[107] = shifted_input7;
      input_sum_parallel[108] = 0;
      input_sum_parallel[109] = shifted_input7;
      input_sum_parallel[110] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[111] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[112] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[113] = shifted_input7;
      input_sum_parallel[114] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[115] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[116] = shifted_input7;
      input_sum_parallel[117] = shifted_input7;
      input_sum_parallel[118] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[119] = shifted_input7;
      input_sum_parallel[120] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[121] = shifted_input7;
      input_sum_parallel[122] = shifted_input7;
      input_sum_parallel[123] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[124] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[125] = shifted_input7;
      input_sum_parallel[126] = shifted_input7;
      input_sum_parallel[127] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[128] = shifted_input7;
      input_sum_parallel[129] = shifted_input7;
      input_sum_parallel[130] = shifted_input7;
      input_sum_parallel[131] = shifted_input7;
      input_sum_parallel[132] = shifted_input7;
      input_sum_parallel[133] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[134] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[135] = shifted_input7;
      input_sum_parallel[136] = shifted_input7;
      input_sum_parallel[137] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[138] = 0;
      input_sum_parallel[139] = shifted_input7;
      input_sum_parallel[140] = shifted_input7;
      input_sum_parallel[141] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[142] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[143] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[144] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[145] = shifted_input7;
      input_sum_parallel[146] = shifted_input7;
      input_sum_parallel[147] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[148] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[149] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[150] = shifted_input7;
      input_sum_parallel[151] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[152] = shifted_input7;
      input_sum_parallel[153] = 0;
      input_sum_parallel[154] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[155] = shifted_input7;
      input_sum_parallel[156] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[157] = shifted_input7;
      input_sum_parallel[158] = shifted_input7;
      input_sum_parallel[159] = shifted_input7;
      input_sum_parallel[160] = shifted_input7;
      input_sum_parallel[161] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[162] = 0;
      input_sum_parallel[163] = shifted_input7;
      input_sum_parallel[164] = 0;
      input_sum_parallel[165] = shifted_input7;
      input_sum_parallel[166] = shifted_input7;
      input_sum_parallel[167] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[168] = shifted_input7;
      input_sum_parallel[169] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[170] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[171] = shifted_input7;
      input_sum_parallel[172] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[173] = shifted_input7;
      input_sum_parallel[174] = shifted_input7;
      input_sum_parallel[175] = 0;
      input_sum_parallel[176] = 0;
      input_sum_parallel[177] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[178] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[179] = shifted_input7;
      input_sum_parallel[180] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[181] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[182] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[183] = 0;
      input_sum_parallel[184] = shifted_input7;
      input_sum_parallel[185] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[186] = shifted_input7;
      input_sum_parallel[187] = shifted_input7;
      input_sum_parallel[188] = shifted_input7;
      input_sum_parallel[189] = shifted_input7;
      input_sum_parallel[190] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[191] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[192] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[193] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
      input_sum_parallel[194] = shifted_input7;
      input_sum_parallel[195] = shifted_input7;
      input_sum_parallel[196] = shifted_input7;
      input_sum_parallel[197] = shifted_input7;
      input_sum_parallel[198] = shifted_input7;
      input_sum_parallel[199] = shifted_input0 + shifted_input1 + shifted_input2 + shifted_input3 + shifted_input4 + shifted_input5 + shifted_input6;
reservoir_sum_parallel[0] = 32'sd0;
reservoir_sum_parallel[1] = 32'sd0;
reservoir_sum_parallel[2] = 32'sd0;
reservoir_sum_parallel[3] = 32'sd0;
reservoir_sum_parallel[4] = 32'sd0;
reservoir_sum_parallel[5] = 32'sd0;
reservoir_sum_parallel[6] = 32'sd0;
reservoir_sum_parallel[7] = 32'sd0;
reservoir_sum_parallel[8] = 32'sd0;
reservoir_sum_parallel[9] = 32'sd0;
reservoir_sum_parallel[10] = 32'sd0;
reservoir_sum_parallel[11] = 32'sd0;
reservoir_sum_parallel[12] = 32'sd0;
reservoir_sum_parallel[13] = 32'sd0;
reservoir_sum_parallel[14] = 32'sd0;
reservoir_sum_parallel[15] = 32'sd0;
reservoir_sum_parallel[16] = 32'sd0;
reservoir_sum_parallel[17] = 32'sd0;
reservoir_sum_parallel[18] = 32'sd0;
reservoir_sum_parallel[19] = 32'sd0;
reservoir_sum_parallel[20] = 32'sd0;
reservoir_sum_parallel[21] = 32'sd0;
reservoir_sum_parallel[22] = 32'sd0;
reservoir_sum_parallel[23] = 32'sd0;
reservoir_sum_parallel[24] = 32'sd0;
reservoir_sum_parallel[25] = 32'sd0;
reservoir_sum_parallel[26] = 32'sd0;
reservoir_sum_parallel[27] = 32'sd0;
reservoir_sum_parallel[28] = 32'sd0;
reservoir_sum_parallel[29] = 32'sd0;
reservoir_sum_parallel[30] = 32'sd0;
reservoir_sum_parallel[31] = 32'sd0;
reservoir_sum_parallel[32] = 32'sd0;
reservoir_sum_parallel[33] = 32'sd0;
reservoir_sum_parallel[34] = 32'sd0;
reservoir_sum_parallel[35] = 32'sd0;
reservoir_sum_parallel[36] = 32'sd0;
reservoir_sum_parallel[37] = 32'sd0;
reservoir_sum_parallel[38] = 32'sd0;
reservoir_sum_parallel[39] = 32'sd0;
reservoir_sum_parallel[40] = 32'sd0;
reservoir_sum_parallel[41] = 32'sd0;
reservoir_sum_parallel[42] = 32'sd0;
reservoir_sum_parallel[43] = 32'sd0;
reservoir_sum_parallel[44] = 32'sd0;
reservoir_sum_parallel[45] = 32'sd0;
reservoir_sum_parallel[46] = 32'sd0;
reservoir_sum_parallel[47] = 32'sd0;
reservoir_sum_parallel[48] = 32'sd0;
reservoir_sum_parallel[49] = 32'sd0;
reservoir_sum_parallel[50] = 32'sd0;
reservoir_sum_parallel[51] = 32'sd0;
reservoir_sum_parallel[52] = 32'sd0;
reservoir_sum_parallel[53] = 32'sd0;
reservoir_sum_parallel[54] = 32'sd0;
reservoir_sum_parallel[55] = 32'sd0;
reservoir_sum_parallel[56] = 32'sd0;
reservoir_sum_parallel[57] = 32'sd0;
reservoir_sum_parallel[58] = 32'sd0;
reservoir_sum_parallel[59] = 32'sd0;
reservoir_sum_parallel[60] = 32'sd0;
reservoir_sum_parallel[61] = 32'sd0;
reservoir_sum_parallel[62] = 32'sd0;
reservoir_sum_parallel[63] = 32'sd0;
reservoir_sum_parallel[64] = 32'sd0;
reservoir_sum_parallel[65] = 32'sd0;
reservoir_sum_parallel[66] = 32'sd0;
reservoir_sum_parallel[67] = 32'sd0;
reservoir_sum_parallel[68] = 32'sd0;
reservoir_sum_parallel[69] = 32'sd0;
reservoir_sum_parallel[70] = 32'sd0;
reservoir_sum_parallel[71] = 32'sd0;
reservoir_sum_parallel[72] = 32'sd0;
reservoir_sum_parallel[73] = 32'sd0;
reservoir_sum_parallel[74] = 32'sd0;
reservoir_sum_parallel[75] = 32'sd0;
reservoir_sum_parallel[76] = 32'sd0;
reservoir_sum_parallel[77] = 32'sd0;
reservoir_sum_parallel[78] = 32'sd0;
reservoir_sum_parallel[79] = 32'sd0;
reservoir_sum_parallel[80] = 32'sd0;
reservoir_sum_parallel[81] = 32'sd0;
reservoir_sum_parallel[82] = 32'sd0;
reservoir_sum_parallel[83] = 32'sd0;
reservoir_sum_parallel[84] = 32'sd0;
reservoir_sum_parallel[85] = 32'sd0;
reservoir_sum_parallel[86] = 32'sd0;
reservoir_sum_parallel[87] = 32'sd0;
reservoir_sum_parallel[88] = 32'sd0;
reservoir_sum_parallel[89] = 32'sd0;
reservoir_sum_parallel[90] = 32'sd0;
reservoir_sum_parallel[91] = 32'sd0;
reservoir_sum_parallel[92] = 32'sd0;
reservoir_sum_parallel[93] = 32'sd0;
reservoir_sum_parallel[94] = 32'sd0;
reservoir_sum_parallel[95] = 32'sd0;
reservoir_sum_parallel[96] = 32'sd0;
reservoir_sum_parallel[97] = 32'sd0;
reservoir_sum_parallel[98] = 32'sd0;
reservoir_sum_parallel[99] = 32'sd0;
reservoir_sum_parallel[100] = 32'sd0;
reservoir_sum_parallel[101] = 32'sd0;
reservoir_sum_parallel[102] = 32'sd0;
reservoir_sum_parallel[103] = 32'sd0;
reservoir_sum_parallel[104] = 32'sd0;
reservoir_sum_parallel[105] = 32'sd0;
reservoir_sum_parallel[106] = 32'sd0;
reservoir_sum_parallel[107] = 32'sd0;
reservoir_sum_parallel[108] = 32'sd0;
reservoir_sum_parallel[109] = 32'sd0;
reservoir_sum_parallel[110] = 32'sd0;
reservoir_sum_parallel[111] = 32'sd0;
reservoir_sum_parallel[112] = 32'sd0;
reservoir_sum_parallel[113] = 32'sd0;
reservoir_sum_parallel[114] = 32'sd0;
reservoir_sum_parallel[115] = 32'sd0;
reservoir_sum_parallel[116] = 32'sd0;
reservoir_sum_parallel[117] = 32'sd0;
reservoir_sum_parallel[118] = 32'sd0;
reservoir_sum_parallel[119] = 32'sd0;
reservoir_sum_parallel[120] = 32'sd0;
reservoir_sum_parallel[121] = 32'sd0;
reservoir_sum_parallel[122] = 32'sd0;
reservoir_sum_parallel[123] = 32'sd0;
reservoir_sum_parallel[124] = 32'sd0;
reservoir_sum_parallel[125] = 32'sd0;
reservoir_sum_parallel[126] = 32'sd0;
reservoir_sum_parallel[127] = 32'sd0;
reservoir_sum_parallel[128] = 32'sd0;
reservoir_sum_parallel[129] = 32'sd0;
reservoir_sum_parallel[130] = 32'sd0;
reservoir_sum_parallel[131] = 32'sd0;
reservoir_sum_parallel[132] = 32'sd0;
reservoir_sum_parallel[133] = 32'sd0;
reservoir_sum_parallel[134] = 32'sd0;
reservoir_sum_parallel[135] = 32'sd0;
reservoir_sum_parallel[136] = 32'sd0;
reservoir_sum_parallel[137] = 32'sd0;
reservoir_sum_parallel[138] = 32'sd0;
reservoir_sum_parallel[139] = 32'sd0;
reservoir_sum_parallel[140] = 32'sd0;
reservoir_sum_parallel[141] = 32'sd0;
reservoir_sum_parallel[142] = 32'sd0;
reservoir_sum_parallel[143] = 32'sd0;
reservoir_sum_parallel[144] = 32'sd0;
reservoir_sum_parallel[145] = 32'sd0;
reservoir_sum_parallel[146] = 32'sd0;
reservoir_sum_parallel[147] = 32'sd0;
reservoir_sum_parallel[148] = 32'sd0;
reservoir_sum_parallel[149] = 32'sd0;
reservoir_sum_parallel[150] = 32'sd0;
reservoir_sum_parallel[151] = 32'sd0;
reservoir_sum_parallel[152] = 32'sd0;
reservoir_sum_parallel[153] = 32'sd0;
reservoir_sum_parallel[154] = 32'sd0;
reservoir_sum_parallel[155] = 32'sd0;
reservoir_sum_parallel[156] = 32'sd0;
reservoir_sum_parallel[157] = 32'sd0;
reservoir_sum_parallel[158] = 32'sd0;
reservoir_sum_parallel[159] = 32'sd0;
reservoir_sum_parallel[160] = 32'sd0;
reservoir_sum_parallel[161] = 32'sd0;
reservoir_sum_parallel[162] = 32'sd0;
reservoir_sum_parallel[163] = 32'sd0;
reservoir_sum_parallel[164] = 32'sd0;
reservoir_sum_parallel[165] = 32'sd0;
reservoir_sum_parallel[166] = 32'sd0;
reservoir_sum_parallel[167] = 32'sd0;
reservoir_sum_parallel[168] = 32'sd0;
reservoir_sum_parallel[169] = 32'sd0;
reservoir_sum_parallel[170] = 32'sd0;
reservoir_sum_parallel[171] = 32'sd0;
reservoir_sum_parallel[172] = 32'sd0;
reservoir_sum_parallel[173] = 32'sd0;
reservoir_sum_parallel[174] = 32'sd0;
reservoir_sum_parallel[175] = 32'sd0;
reservoir_sum_parallel[176] = 32'sd0;
reservoir_sum_parallel[177] = 32'sd0;
reservoir_sum_parallel[178] = 32'sd0;
reservoir_sum_parallel[179] = 32'sd0;
reservoir_sum_parallel[180] = 32'sd0;
reservoir_sum_parallel[181] = 32'sd0;
reservoir_sum_parallel[182] = 32'sd0;
reservoir_sum_parallel[183] = 32'sd0;
reservoir_sum_parallel[184] = 32'sd0;
reservoir_sum_parallel[185] = 32'sd0;
reservoir_sum_parallel[186] = 32'sd0;
reservoir_sum_parallel[187] = 32'sd0;
reservoir_sum_parallel[188] = 32'sd0;
reservoir_sum_parallel[189] = 32'sd0;
reservoir_sum_parallel[190] = 32'sd0;
reservoir_sum_parallel[191] = 32'sd0;
reservoir_sum_parallel[192] = 32'sd0;
reservoir_sum_parallel[193] = 32'sd0;
reservoir_sum_parallel[194] = 32'sd0;
reservoir_sum_parallel[195] = 32'sd0;
reservoir_sum_parallel[196] = 32'sd0;
reservoir_sum_parallel[197] = 32'sd0;
reservoir_sum_parallel[198] = 32'sd0;
reservoir_sum_parallel[199] = 32'sd0;
      reservoir_sum_parallel[0] = (shifted_state0_19_0 + shifted_state0_19_3 + shifted_state0_19_4 + shifted_state0_19_6 + shifted_state0_19_7 + shifted_state0_40_0 + shifted_state0_40_1 + shifted_state0_40_2 + shifted_state0_40_3 + shifted_state0_40_4 + shifted_state0_47_0 + shifted_state0_47_1 + shifted_state0_47_2 + shifted_state0_47_4 + shifted_state0_47_5 + shifted_state0_47_6 + shifted_state0_47_7 + shifted_state0_59_0 + shifted_state0_59_4 + shifted_state0_59_5 + shifted_state0_59_7 + shifted_state0_63_1 + shifted_state0_63_3 + shifted_state0_63_4 + shifted_state0_87_3 + shifted_state0_87_5 + shifted_state0_87_6 + shifted_state0_87_7 + shifted_state0_115_4 + shifted_state0_115_5 + shifted_state0_115_6 + shifted_state0_115_7 + shifted_state0_117_0 + shifted_state0_117_1 + shifted_state0_117_2 + shifted_state0_117_3 + shifted_state0_117_4 + shifted_state0_117_5 + shifted_state0_117_6 + shifted_state0_117_7 + shifted_state0_124_0 + shifted_state0_124_1 + shifted_state0_124_5 + shifted_state0_153_1 + shifted_state0_153_2 + shifted_state0_153_3 + shifted_state0_153_4 + shifted_state0_158_1 + shifted_state0_158_2 + shifted_state0_158_5 + shifted_state0_171_0 + shifted_state0_172_1 + shifted_state0_174_1 + shifted_state0_174_2 + shifted_state0_174_4 + shifted_state0_174_5 + shifted_state0_174_6 + shifted_state0_174_7 + shifted_state0_176_1 + shifted_state0_176_2 + shifted_state0_176_5 + shifted_state0_176_6 + shifted_state0_176_7 + shifted_state0_182_3 + shifted_state0_191_1 + shifted_state0_191_2 + shifted_state0_191_3 + shifted_state0_191_4 + shifted_state0_191_5 + shifted_state0_191_6 + shifted_state0_191_7 + shifted_state0_196_3 + shifted_state0_196_6);
      reservoir_sum_parallel[1] = (shifted_state1_4_0 + shifted_state1_4_1 + shifted_state1_4_4 + shifted_state1_4_5 + shifted_state1_4_6 + shifted_state1_4_7 + shifted_state1_10_0 + shifted_state1_10_5 + shifted_state1_12_1 + shifted_state1_12_4 + shifted_state1_14_0 + shifted_state1_14_1 + shifted_state1_14_3 + shifted_state1_14_4 + shifted_state1_14_5 + shifted_state1_14_6 + shifted_state1_14_7 + shifted_state1_42_0 + shifted_state1_42_1 + shifted_state1_42_3 + shifted_state1_42_4 + shifted_state1_57_0 + shifted_state1_57_3 + shifted_state1_57_4 + shifted_state1_57_5 + shifted_state1_57_6 + shifted_state1_57_7 + shifted_state1_78_2 + shifted_state1_78_5 + shifted_state1_83_0 + shifted_state1_83_1 + shifted_state1_83_3 + shifted_state1_91_0 + shifted_state1_91_1 + shifted_state1_91_6 + shifted_state1_91_7 + shifted_state1_93_0 + shifted_state1_93_1 + shifted_state1_93_2 + shifted_state1_93_3 + shifted_state1_93_4 + shifted_state1_108_0 + shifted_state1_108_3 + shifted_state1_114_0 + shifted_state1_114_1 + shifted_state1_114_3 + shifted_state1_119_1 + shifted_state1_119_2 + shifted_state1_119_3 + shifted_state1_127_0 + shifted_state1_127_2 + shifted_state1_127_3 + shifted_state1_127_4 + shifted_state1_127_5 + shifted_state1_127_6 + shifted_state1_127_7 + shifted_state1_131_1 + shifted_state1_131_2 + shifted_state1_131_4 + shifted_state1_131_5 + shifted_state1_131_6 + shifted_state1_131_7 + shifted_state1_154_1 + shifted_state1_154_2 + shifted_state1_154_3 + shifted_state1_154_5 + shifted_state1_154_6 + shifted_state1_154_7 + shifted_state1_156_2 + shifted_state1_156_3 + shifted_state1_156_5 + shifted_state1_156_6 + shifted_state1_156_7 + shifted_state1_165_1 + shifted_state1_165_3 + shifted_state1_189_0 + shifted_state1_189_4 + shifted_state1_193_0 + shifted_state1_193_1 + shifted_state1_193_2 + shifted_state1_193_4 + shifted_state1_198_0 + shifted_state1_198_3);
      reservoir_sum_parallel[2] = (shifted_state2_17_1 + shifted_state2_17_2 + shifted_state2_17_4 + shifted_state2_17_5 + shifted_state2_17_6 + shifted_state2_17_7 + shifted_state2_35_2 + shifted_state2_35_3 + shifted_state2_35_4 + shifted_state2_35_6 + shifted_state2_35_7 + shifted_state2_73_0 + shifted_state2_73_1 + shifted_state2_73_4 + shifted_state2_77_1 + shifted_state2_77_2 + shifted_state2_77_4 + shifted_state2_77_5 + shifted_state2_82_2 + shifted_state2_82_3 + shifted_state2_82_5 + shifted_state2_82_6 + shifted_state2_82_7 + shifted_state2_132_3 + shifted_state2_132_5 + shifted_state2_140_0 + shifted_state2_140_4 + shifted_state2_140_6 + shifted_state2_140_7 + shifted_state2_151_0 + shifted_state2_151_4 + shifted_state2_151_5 + shifted_state2_170_0 + shifted_state2_170_1 + shifted_state2_170_2 + shifted_state2_170_4 + shifted_state2_172_0 + shifted_state2_172_1 + shifted_state2_172_2 + shifted_state2_172_3 + shifted_state2_172_4 + shifted_state2_172_5 + shifted_state2_172_6 + shifted_state2_172_7 + shifted_state2_182_0 + shifted_state2_182_3 + shifted_state2_182_4);
      reservoir_sum_parallel[3] = (shifted_state3_15_1 + shifted_state3_15_6 + shifted_state3_15_7 + shifted_state3_31_4 + shifted_state3_31_5 + shifted_state3_31_6 + shifted_state3_31_7 + shifted_state3_36_0 + shifted_state3_36_2 + shifted_state3_36_3 + shifted_state3_36_4 + shifted_state3_36_6 + shifted_state3_36_7 + shifted_state3_41_0 + shifted_state3_41_2 + shifted_state3_41_3 + shifted_state3_41_4 + shifted_state3_41_5 + shifted_state3_41_6 + shifted_state3_41_7 + shifted_state3_44_0 + shifted_state3_44_1 + shifted_state3_44_3 + shifted_state3_44_6 + shifted_state3_44_7 + shifted_state3_66_0 + shifted_state3_66_3 + shifted_state3_66_5 + shifted_state3_66_6 + shifted_state3_66_7 + shifted_state3_82_0 + shifted_state3_82_1 + shifted_state3_82_4 + shifted_state3_82_5 + shifted_state3_82_6 + shifted_state3_82_7 + shifted_state3_96_0 + shifted_state3_96_1 + shifted_state3_96_2 + shifted_state3_96_3 + shifted_state3_96_5 + shifted_state3_96_6 + shifted_state3_96_7 + shifted_state3_104_0 + shifted_state3_104_1 + shifted_state3_104_4 + shifted_state3_111_2 + shifted_state3_131_1 + shifted_state3_131_3 + shifted_state3_149_5 + shifted_state3_149_6 + shifted_state3_149_7 + shifted_state3_166_1 + shifted_state3_166_2 + shifted_state3_166_3 + shifted_state3_166_6 + shifted_state3_166_7 + shifted_state3_186_0 + shifted_state3_186_2 + shifted_state3_186_4 + shifted_state3_190_0 + shifted_state3_190_2 + shifted_state3_190_4 + shifted_state3_190_5 + shifted_state3_191_0 + shifted_state3_191_2);
      reservoir_sum_parallel[4] = (shifted_state4_4_1 + shifted_state4_4_2 + shifted_state4_4_3 + shifted_state4_4_4 + shifted_state4_4_5 + shifted_state4_4_6 + shifted_state4_4_7 + shifted_state4_34_4 + shifted_state4_34_6 + shifted_state4_34_7 + shifted_state4_41_0 + shifted_state4_41_1 + shifted_state4_41_5 + shifted_state4_51_1 + shifted_state4_51_3 + shifted_state4_51_4 + shifted_state4_51_5 + shifted_state4_58_0 + shifted_state4_58_1 + shifted_state4_58_3 + shifted_state4_58_4 + shifted_state4_58_5 + shifted_state4_58_6 + shifted_state4_58_7 + shifted_state4_66_4 + shifted_state4_66_5 + shifted_state4_72_4 + shifted_state4_76_4 + shifted_state4_76_5 + shifted_state4_76_6 + shifted_state4_76_7 + shifted_state4_79_0 + shifted_state4_79_2 + shifted_state4_85_0 + shifted_state4_85_3 + shifted_state4_93_3 + shifted_state4_96_0 + shifted_state4_96_2 + shifted_state4_96_5 + shifted_state4_104_2 + shifted_state4_104_4 + shifted_state4_104_5 + shifted_state4_105_1 + shifted_state4_105_2 + shifted_state4_105_5 + shifted_state4_105_6 + shifted_state4_105_7 + shifted_state4_119_3 + shifted_state4_119_4 + shifted_state4_119_5 + shifted_state4_119_6 + shifted_state4_119_7 + shifted_state4_139_4 + shifted_state4_139_5 + shifted_state4_139_6 + shifted_state4_139_7 + shifted_state4_163_0 + shifted_state4_163_2 + shifted_state4_163_4 + shifted_state4_165_1 + shifted_state4_165_3 + shifted_state4_183_0 + shifted_state4_183_1 + shifted_state4_183_2 + shifted_state4_183_3 + shifted_state4_183_4 + shifted_state4_183_5 + shifted_state4_183_7 + shifted_state4_191_0 + shifted_state4_191_1 + shifted_state4_191_2 + shifted_state4_191_4 + shifted_state4_192_0 + shifted_state4_193_0 + shifted_state4_193_2 + shifted_state4_193_3 + shifted_state4_197_0 + shifted_state4_197_1 + shifted_state4_197_4 + shifted_state4_197_6 + shifted_state4_199_0 + shifted_state4_199_2 + shifted_state4_199_3 + shifted_state4_199_5 + shifted_state4_199_6 + shifted_state4_199_7);
      reservoir_sum_parallel[5] = (shifted_state5_12_0 + shifted_state5_12_2 + shifted_state5_12_4 + shifted_state5_97_1 + shifted_state5_97_4 + shifted_state5_126_5 + shifted_state5_128_6 + shifted_state5_128_7 + shifted_state5_135_0 + shifted_state5_135_1 + shifted_state5_135_3 + shifted_state5_135_5 + shifted_state5_143_0 + shifted_state5_143_1 + shifted_state5_143_2 + shifted_state5_145_1 + shifted_state5_145_2 + shifted_state5_145_3 + shifted_state5_145_4 + shifted_state5_145_5 + shifted_state5_145_6 + shifted_state5_145_7 + shifted_state5_150_3 + shifted_state5_150_5 + shifted_state5_150_6 + shifted_state5_150_7 + shifted_state5_162_1 + shifted_state5_162_2 + shifted_state5_162_5 + shifted_state5_162_6 + shifted_state5_162_7 + shifted_state5_166_3 + shifted_state5_166_4 + shifted_state5_166_5 + shifted_state5_166_6 + shifted_state5_166_7 + shifted_state5_167_1 + shifted_state5_167_3 + shifted_state5_167_4 + shifted_state5_199_0 + shifted_state5_199_1 + shifted_state5_199_2 + shifted_state5_199_6 + shifted_state5_199_7);
      reservoir_sum_parallel[6] = (shifted_state6_3_3 + shifted_state6_3_5 + shifted_state6_12_0 + shifted_state6_12_1 + shifted_state6_12_2 + shifted_state6_28_3 + shifted_state6_28_4 + shifted_state6_28_5 + shifted_state6_28_6 + shifted_state6_28_7 + shifted_state6_64_0 + shifted_state6_64_3 + shifted_state6_64_4 + shifted_state6_69_1 + shifted_state6_69_2 + shifted_state6_69_3 + shifted_state6_69_4 + shifted_state6_88_0 + shifted_state6_88_1 + shifted_state6_88_5 + shifted_state6_106_2 + shifted_state6_106_3 + shifted_state6_106_4 + shifted_state6_112_2 + shifted_state6_112_3 + shifted_state6_112_4 + shifted_state6_112_5 + shifted_state6_112_6 + shifted_state6_112_7 + shifted_state6_136_3 + shifted_state6_136_5 + shifted_state6_136_6 + shifted_state6_136_7 + shifted_state6_147_2 + shifted_state6_147_3 + shifted_state6_150_0 + shifted_state6_150_5 + shifted_state6_158_1 + shifted_state6_158_2 + shifted_state6_158_5 + shifted_state6_158_6 + shifted_state6_158_7 + shifted_state6_168_4 + shifted_state6_168_5 + shifted_state6_168_6 + shifted_state6_168_7 + shifted_state6_181_1 + shifted_state6_181_4 + shifted_state6_182_4 + shifted_state6_182_5 + shifted_state6_182_6 + shifted_state6_182_7 + shifted_state6_192_0 + shifted_state6_192_1 + shifted_state6_192_3 + shifted_state6_192_4 + shifted_state6_192_5 + shifted_state6_192_6 + shifted_state6_192_7);
      reservoir_sum_parallel[7] = (shifted_state7_7_2 + shifted_state7_7_3 + shifted_state7_16_0 + shifted_state7_16_3 + shifted_state7_16_4 + shifted_state7_16_5 + shifted_state7_16_6 + shifted_state7_16_7 + shifted_state7_20_1 + shifted_state7_32_0 + shifted_state7_32_1 + shifted_state7_32_2 + shifted_state7_32_3 + shifted_state7_32_5 + shifted_state7_32_6 + shifted_state7_32_7 + shifted_state7_40_3 + shifted_state7_80_0 + shifted_state7_80_1 + shifted_state7_80_3 + shifted_state7_80_4 + shifted_state7_80_5 + shifted_state7_80_6 + shifted_state7_80_7 + shifted_state7_84_7 + shifted_state7_86_0 + shifted_state7_86_1 + shifted_state7_86_2 + shifted_state7_86_3 + shifted_state7_86_4 + shifted_state7_86_5 + shifted_state7_86_6 + shifted_state7_86_7 + shifted_state7_94_1 + shifted_state7_94_2 + shifted_state7_94_3 + shifted_state7_94_4 + shifted_state7_94_5 + shifted_state7_94_6 + shifted_state7_94_7 + shifted_state7_104_4 + shifted_state7_108_0 + shifted_state7_108_2 + shifted_state7_108_5 + shifted_state7_128_0 + shifted_state7_128_2 + shifted_state7_128_3 + shifted_state7_128_5 + shifted_state7_128_6 + shifted_state7_128_7 + shifted_state7_137_1 + shifted_state7_137_3 + shifted_state7_137_4 + shifted_state7_137_6 + shifted_state7_137_7 + shifted_state7_171_1 + shifted_state7_171_2 + shifted_state7_171_5 + shifted_state7_183_0 + shifted_state7_183_1 + shifted_state7_183_2 + shifted_state7_183_4 + shifted_state7_187_4 + shifted_state7_187_5);
      reservoir_sum_parallel[8] = (shifted_state8_3_0 + shifted_state8_3_2 + shifted_state8_3_4 + shifted_state8_3_6 + shifted_state8_3_7 + shifted_state8_24_0 + shifted_state8_24_1 + shifted_state8_24_2 + shifted_state8_36_0 + shifted_state8_36_1 + shifted_state8_36_5 + shifted_state8_45_1 + shifted_state8_45_2 + shifted_state8_45_3 + shifted_state8_45_4 + shifted_state8_53_0 + shifted_state8_53_3 + shifted_state8_54_0 + shifted_state8_54_1 + shifted_state8_54_2 + shifted_state8_55_0 + shifted_state8_55_1 + shifted_state8_55_3 + shifted_state8_55_5 + shifted_state8_55_6 + shifted_state8_55_7 + shifted_state8_56_1 + shifted_state8_56_2 + shifted_state8_56_3 + shifted_state8_56_4 + shifted_state8_61_0 + shifted_state8_61_1 + shifted_state8_61_2 + shifted_state8_61_4 + shifted_state8_79_0 + shifted_state8_79_2 + shifted_state8_79_3 + shifted_state8_79_6 + shifted_state8_79_7 + shifted_state8_88_0 + shifted_state8_93_0 + shifted_state8_93_1 + shifted_state8_93_2 + shifted_state8_93_3 + shifted_state8_93_5 + shifted_state8_93_6 + shifted_state8_93_7 + shifted_state8_96_1 + shifted_state8_96_2 + shifted_state8_96_3 + shifted_state8_114_3 + shifted_state8_114_5 + shifted_state8_114_6 + shifted_state8_114_7 + shifted_state8_125_0 + shifted_state8_125_2 + shifted_state8_125_3 + shifted_state8_125_6 + shifted_state8_125_7 + shifted_state8_131_0 + shifted_state8_131_1 + shifted_state8_131_2 + shifted_state8_131_3 + shifted_state8_131_6 + shifted_state8_131_7 + shifted_state8_136_0 + shifted_state8_136_3 + shifted_state8_136_4 + shifted_state8_149_0 + shifted_state8_149_2 + shifted_state8_149_3 + shifted_state8_173_0 + shifted_state8_173_1 + shifted_state8_173_2 + shifted_state8_173_3 + shifted_state8_173_5 + shifted_state8_173_6 + shifted_state8_173_7 + shifted_state8_180_0 + shifted_state8_180_1 + shifted_state8_180_3 + shifted_state8_187_0 + shifted_state8_187_5 + shifted_state8_187_6 + shifted_state8_187_7);
      reservoir_sum_parallel[9] = (shifted_state9_22_2 + shifted_state9_22_4 + shifted_state9_22_6 + shifted_state9_22_7 + shifted_state9_23_1 + shifted_state9_23_2 + shifted_state9_31_0 + shifted_state9_31_1 + shifted_state9_31_3 + shifted_state9_31_5 + shifted_state9_31_6 + shifted_state9_31_7 + shifted_state9_52_0 + shifted_state9_52_1 + shifted_state9_52_3 + shifted_state9_52_4 + shifted_state9_59_2 + shifted_state9_59_3 + shifted_state9_69_3 + shifted_state9_69_4 + shifted_state9_71_0 + shifted_state9_71_1 + shifted_state9_71_2 + shifted_state9_71_3 + shifted_state9_71_4 + shifted_state9_82_3 + shifted_state9_86_0 + shifted_state9_86_1 + shifted_state9_86_3 + shifted_state9_86_5 + shifted_state9_86_6 + shifted_state9_86_7 + shifted_state9_95_0 + shifted_state9_95_3 + shifted_state9_95_5 + shifted_state9_95_6 + shifted_state9_95_7 + shifted_state9_105_0 + shifted_state9_105_1 + shifted_state9_105_2 + shifted_state9_105_4 + shifted_state9_107_1 + shifted_state9_107_4 + shifted_state9_107_6 + shifted_state9_107_7 + shifted_state9_137_0 + shifted_state9_137_1 + shifted_state9_137_2 + shifted_state9_139_1 + shifted_state9_139_4 + shifted_state9_141_0 + shifted_state9_141_2 + shifted_state9_141_3 + shifted_state9_141_5 + shifted_state9_141_6 + shifted_state9_141_7 + shifted_state9_163_1 + shifted_state9_163_2 + shifted_state9_163_5 + shifted_state9_163_6 + shifted_state9_163_7 + shifted_state9_165_1 + shifted_state9_165_2 + shifted_state9_165_3 + shifted_state9_170_1 + shifted_state9_170_2 + shifted_state9_170_3 + shifted_state9_175_1 + shifted_state9_175_3 + shifted_state9_175_4 + shifted_state9_175_6 + shifted_state9_175_7 + shifted_state9_188_1 + shifted_state9_188_4 + shifted_state9_190_0 + shifted_state9_190_1 + shifted_state9_190_3 + shifted_state9_190_5 + shifted_state9_190_6 + shifted_state9_190_7);
      reservoir_sum_parallel[10] = (shifted_state10_17_1 + shifted_state10_17_2 + shifted_state10_17_3 + shifted_state10_22_0 + shifted_state10_22_2 + shifted_state10_22_4 + shifted_state10_22_5 + shifted_state10_22_6 + shifted_state10_22_7 + shifted_state10_40_1 + shifted_state10_40_3 + shifted_state10_48_0 + shifted_state10_48_3 + shifted_state10_56_0 + shifted_state10_56_1 + shifted_state10_56_2 + shifted_state10_73_0 + shifted_state10_73_3 + shifted_state10_73_6 + shifted_state10_73_7 + shifted_state10_74_2 + shifted_state10_74_3 + shifted_state10_74_5 + shifted_state10_74_6 + shifted_state10_74_7 + shifted_state10_78_3 + shifted_state10_78_6 + shifted_state10_78_7 + shifted_state10_106_0 + shifted_state10_106_1 + shifted_state10_106_2 + shifted_state10_106_3 + shifted_state10_121_0 + shifted_state10_121_2 + shifted_state10_121_4 + shifted_state10_121_5 + shifted_state10_121_6 + shifted_state10_121_7 + shifted_state10_131_0 + shifted_state10_131_2 + shifted_state10_131_4 + shifted_state10_131_5 + shifted_state10_131_6 + shifted_state10_131_7 + shifted_state10_132_1 + shifted_state10_132_3 + shifted_state10_132_4 + shifted_state10_132_5 + shifted_state10_132_6 + shifted_state10_132_7 + shifted_state10_133_0 + shifted_state10_133_4 + shifted_state10_165_0 + shifted_state10_165_1 + shifted_state10_165_2 + shifted_state10_165_3 + shifted_state10_165_4 + shifted_state10_170_0 + shifted_state10_170_3 + shifted_state10_176_0 + shifted_state10_176_1 + shifted_state10_176_4 + shifted_state10_176_5 + shifted_state10_176_6 + shifted_state10_176_7 + shifted_state10_177_0 + shifted_state10_177_4 + shifted_state10_179_2 + shifted_state10_179_3 + shifted_state10_179_5 + shifted_state10_179_6 + shifted_state10_179_7 + shifted_state10_180_0 + shifted_state10_180_2 + shifted_state10_180_4 + shifted_state10_180_5 + shifted_state10_180_6 + shifted_state10_180_7 + shifted_state10_185_0 + shifted_state10_185_1 + shifted_state10_185_3 + shifted_state10_185_4 + shifted_state10_186_0 + shifted_state10_186_1 + shifted_state10_186_3 + shifted_state10_186_6 + shifted_state10_186_7);
      reservoir_sum_parallel[11] = (shifted_state11_26_1 + shifted_state11_26_2 + shifted_state11_26_3 + shifted_state11_26_5 + shifted_state11_26_6 + shifted_state11_26_7 + shifted_state11_31_2 + shifted_state11_31_4 + shifted_state11_31_5 + shifted_state11_31_6 + shifted_state11_31_7 + shifted_state11_33_0 + shifted_state11_33_1 + shifted_state11_33_2 + shifted_state11_33_3 + shifted_state11_33_4 + shifted_state11_33_5 + shifted_state11_33_6 + shifted_state11_33_7 + shifted_state11_34_0 + shifted_state11_34_2 + shifted_state11_34_3 + shifted_state11_34_5 + shifted_state11_40_0 + shifted_state11_40_1 + shifted_state11_40_6 + shifted_state11_58_3 + shifted_state11_58_4 + shifted_state11_58_6 + shifted_state11_58_7 + shifted_state11_100_1 + shifted_state11_111_0 + shifted_state11_111_2 + shifted_state11_111_6 + shifted_state11_111_7 + shifted_state11_123_0 + shifted_state11_123_2 + shifted_state11_123_4 + shifted_state11_123_5 + shifted_state11_123_6 + shifted_state11_123_7 + shifted_state11_130_0 + shifted_state11_130_2 + shifted_state11_130_3 + shifted_state11_130_4 + shifted_state11_130_5 + shifted_state11_130_6 + shifted_state11_130_7 + shifted_state11_132_0 + shifted_state11_132_2 + shifted_state11_132_3 + shifted_state11_132_5 + shifted_state11_132_6 + shifted_state11_132_7 + shifted_state11_135_0 + shifted_state11_135_4 + shifted_state11_135_6 + shifted_state11_135_7 + shifted_state11_139_4 + shifted_state11_143_3 + shifted_state11_143_5 + shifted_state11_143_6 + shifted_state11_143_7 + shifted_state11_147_0 + shifted_state11_147_2 + shifted_state11_147_5 + shifted_state11_147_6 + shifted_state11_147_7 + shifted_state11_150_0 + shifted_state11_150_2 + shifted_state11_150_3 + shifted_state11_151_3 + shifted_state11_151_5 + shifted_state11_151_6 + shifted_state11_151_7 + shifted_state11_158_2 + shifted_state11_158_4 + shifted_state11_158_5 + shifted_state11_158_6 + shifted_state11_158_7);
      reservoir_sum_parallel[12] = (shifted_state12_6_0 + shifted_state12_6_1 + shifted_state12_6_5 + shifted_state12_6_6 + shifted_state12_6_7 + shifted_state12_7_0 + shifted_state12_7_1 + shifted_state12_7_2 + shifted_state12_7_4 + shifted_state12_28_0 + shifted_state12_28_3 + shifted_state12_28_4 + shifted_state12_54_1 + shifted_state12_54_2 + shifted_state12_54_3 + shifted_state12_54_4 + shifted_state12_54_5 + shifted_state12_54_6 + shifted_state12_54_7 + shifted_state12_63_1 + shifted_state12_63_2 + shifted_state12_63_3 + shifted_state12_75_0 + shifted_state12_75_1 + shifted_state12_75_2 + shifted_state12_75_3 + shifted_state12_75_5 + shifted_state12_82_0 + shifted_state12_82_1 + shifted_state12_82_2 + shifted_state12_82_4 + shifted_state12_82_5 + shifted_state12_82_6 + shifted_state12_82_7 + shifted_state12_86_1 + shifted_state12_86_2 + shifted_state12_86_5 + shifted_state12_86_6 + shifted_state12_86_7 + shifted_state12_125_0 + shifted_state12_125_4 + shifted_state12_125_5 + shifted_state12_125_6 + shifted_state12_125_7 + shifted_state12_130_3 + shifted_state12_130_4 + shifted_state12_130_5 + shifted_state12_130_6 + shifted_state12_130_7 + shifted_state12_144_0 + shifted_state12_144_2 + shifted_state12_144_3 + shifted_state12_144_5 + shifted_state12_144_6 + shifted_state12_144_7 + shifted_state12_150_0 + shifted_state12_150_1 + shifted_state12_150_2 + shifted_state12_150_4 + shifted_state12_150_5 + shifted_state12_150_6 + shifted_state12_150_7 + shifted_state12_165_0 + shifted_state12_165_2 + shifted_state12_165_3 + shifted_state12_165_4 + shifted_state12_165_5 + shifted_state12_165_6 + shifted_state12_165_7 + shifted_state12_169_1 + shifted_state12_169_5 + shifted_state12_175_1 + shifted_state12_175_2 + shifted_state12_175_3 + shifted_state12_175_4 + shifted_state12_175_5 + shifted_state12_175_6 + shifted_state12_175_7 + shifted_state12_180_4 + shifted_state12_180_6 + shifted_state12_180_7 + shifted_state12_182_0 + shifted_state12_182_3 + shifted_state12_187_2 + shifted_state12_187_3 + shifted_state12_192_1 + shifted_state12_192_2 + shifted_state12_192_4 + shifted_state12_192_5 + shifted_state12_192_6 + shifted_state12_192_7 + shifted_state12_195_0 + shifted_state12_195_1 + shifted_state12_195_2 + shifted_state12_195_4 + shifted_state12_195_5 + shifted_state12_195_6 + shifted_state12_195_7 + shifted_state12_197_0 + shifted_state12_197_2 + shifted_state12_197_5 + shifted_state12_199_0 + shifted_state12_199_1 + shifted_state12_199_2 + shifted_state12_199_3 + shifted_state12_199_4 + shifted_state12_199_5 + shifted_state12_199_6 + shifted_state12_199_7);
      reservoir_sum_parallel[13] = (shifted_state13_0_0 + shifted_state13_0_1 + shifted_state13_0_4 + shifted_state13_0_5 + shifted_state13_0_6 + shifted_state13_0_7 + shifted_state13_11_0 + shifted_state13_11_1 + shifted_state13_11_4 + shifted_state13_11_5 + shifted_state13_11_6 + shifted_state13_11_7 + shifted_state13_26_2 + shifted_state13_26_3 + shifted_state13_26_6 + shifted_state13_26_7 + shifted_state13_27_1 + shifted_state13_27_2 + shifted_state13_27_3 + shifted_state13_27_4 + shifted_state13_27_5 + shifted_state13_27_6 + shifted_state13_27_7 + shifted_state13_30_0 + shifted_state13_30_1 + shifted_state13_30_3 + shifted_state13_30_4 + shifted_state13_38_1 + shifted_state13_38_2 + shifted_state13_38_3 + shifted_state13_57_2 + shifted_state13_57_3 + shifted_state13_57_5 + shifted_state13_57_6 + shifted_state13_57_7 + shifted_state13_79_2 + shifted_state13_79_3 + shifted_state13_79_4 + shifted_state13_79_5 + shifted_state13_79_6 + shifted_state13_79_7 + shifted_state13_95_1 + shifted_state13_95_3 + shifted_state13_95_4 + shifted_state13_95_5 + shifted_state13_95_6 + shifted_state13_95_7 + shifted_state13_100_2 + shifted_state13_100_3 + shifted_state13_100_4 + shifted_state13_100_5 + shifted_state13_100_7 + shifted_state13_105_1 + shifted_state13_105_2 + shifted_state13_105_3 + shifted_state13_105_4 + shifted_state13_105_5 + shifted_state13_105_6 + shifted_state13_105_7 + shifted_state13_113_0 + shifted_state13_113_1 + shifted_state13_113_2 + shifted_state13_113_3 + shifted_state13_113_5 + shifted_state13_130_3 + shifted_state13_141_0 + shifted_state13_141_2 + shifted_state13_141_4 + shifted_state13_145_3 + shifted_state13_145_4 + shifted_state13_145_5 + shifted_state13_145_6 + shifted_state13_145_7 + shifted_state13_166_0 + shifted_state13_166_5 + shifted_state13_166_6 + shifted_state13_166_7);
      reservoir_sum_parallel[14] = (shifted_state14_8_4 + shifted_state14_20_0 + shifted_state14_20_3 + shifted_state14_30_2 + shifted_state14_30_5 + shifted_state14_30_6 + shifted_state14_30_7 + shifted_state14_31_0 + shifted_state14_31_3 + shifted_state14_31_4 + shifted_state14_31_5 + shifted_state14_31_7 + shifted_state14_50_1 + shifted_state14_50_3 + shifted_state14_50_5 + shifted_state14_50_6 + shifted_state14_50_7 + shifted_state14_63_3 + shifted_state14_63_4 + shifted_state14_63_6 + shifted_state14_63_7 + shifted_state14_68_0 + shifted_state14_68_1 + shifted_state14_68_3 + shifted_state14_68_6 + shifted_state14_68_7 + shifted_state14_76_0 + shifted_state14_76_4 + shifted_state14_77_3 + shifted_state14_77_4 + shifted_state14_77_5 + shifted_state14_77_6 + shifted_state14_77_7 + shifted_state14_118_1 + shifted_state14_118_6 + shifted_state14_118_7 + shifted_state14_120_0 + shifted_state14_120_1 + shifted_state14_120_3 + shifted_state14_120_4 + shifted_state14_120_5 + shifted_state14_120_6 + shifted_state14_120_7 + shifted_state14_183_0 + shifted_state14_183_1 + shifted_state14_183_6 + shifted_state14_183_7 + shifted_state14_191_0 + shifted_state14_191_3);
      reservoir_sum_parallel[15] = (shifted_state15_0_0 + shifted_state15_0_1 + shifted_state15_0_3 + shifted_state15_0_4 + shifted_state15_0_5 + shifted_state15_0_6 + shifted_state15_0_7 + shifted_state15_4_0 + shifted_state15_4_1 + shifted_state15_4_2 + shifted_state15_4_3 + shifted_state15_5_3 + shifted_state15_5_4 + shifted_state15_5_5 + shifted_state15_5_6 + shifted_state15_5_7 + shifted_state15_7_5 + shifted_state15_26_2 + shifted_state15_26_3 + shifted_state15_26_5 + shifted_state15_48_0 + shifted_state15_48_1 + shifted_state15_48_3 + shifted_state15_53_0 + shifted_state15_53_2 + shifted_state15_53_4 + shifted_state15_99_1 + shifted_state15_99_2 + shifted_state15_99_3 + shifted_state15_99_6 + shifted_state15_99_7 + shifted_state15_111_0 + shifted_state15_111_4 + shifted_state15_111_6 + shifted_state15_111_7 + shifted_state15_114_0 + shifted_state15_114_3 + shifted_state15_114_4 + shifted_state15_114_5 + shifted_state15_114_6 + shifted_state15_114_7 + shifted_state15_119_0 + shifted_state15_119_5 + shifted_state15_121_1 + shifted_state15_121_2 + shifted_state15_121_4 + shifted_state15_121_5 + shifted_state15_121_6 + shifted_state15_121_7 + shifted_state15_153_2 + shifted_state15_153_3 + shifted_state15_153_6 + shifted_state15_153_7 + shifted_state15_154_1 + shifted_state15_157_0 + shifted_state15_157_2 + shifted_state15_157_4 + shifted_state15_157_5 + shifted_state15_157_6 + shifted_state15_157_7 + shifted_state15_184_1 + shifted_state15_184_2 + shifted_state15_184_4 + shifted_state15_193_0 + shifted_state15_193_3 + shifted_state15_193_4 + shifted_state15_193_5 + shifted_state15_193_6 + shifted_state15_193_7 + shifted_state15_197_1 + shifted_state15_197_3 + shifted_state15_197_6 + shifted_state15_197_7 + shifted_state15_199_1);
      reservoir_sum_parallel[16] = (shifted_state16_21_2 + shifted_state16_21_5 + shifted_state16_35_4 + shifted_state16_35_5 + shifted_state16_35_6 + shifted_state16_35_7 + shifted_state16_36_0 + shifted_state16_36_1 + shifted_state16_36_3 + shifted_state16_70_3 + shifted_state16_70_5 + shifted_state16_70_6 + shifted_state16_70_7 + shifted_state16_71_0 + shifted_state16_71_1 + shifted_state16_71_2 + shifted_state16_72_0 + shifted_state16_72_2 + shifted_state16_72_3 + shifted_state16_72_5 + shifted_state16_72_7 + shifted_state16_79_0 + shifted_state16_79_1 + shifted_state16_79_2 + shifted_state16_79_4 + shifted_state16_82_0 + shifted_state16_82_1 + shifted_state16_82_2 + shifted_state16_82_3 + shifted_state16_82_5 + shifted_state16_82_6 + shifted_state16_82_7 + shifted_state16_86_0 + shifted_state16_86_4 + shifted_state16_86_5 + shifted_state16_86_6 + shifted_state16_86_7 + shifted_state16_122_1 + shifted_state16_122_4 + shifted_state16_122_5 + shifted_state16_122_6 + shifted_state16_122_7 + shifted_state16_134_0 + shifted_state16_134_4 + shifted_state16_134_5 + shifted_state16_134_6 + shifted_state16_134_7 + shifted_state16_139_0 + shifted_state16_139_1 + shifted_state16_139_3 + shifted_state16_139_4 + shifted_state16_139_5 + shifted_state16_139_6 + shifted_state16_139_7 + shifted_state16_157_0 + shifted_state16_157_3 + shifted_state16_157_5 + shifted_state16_157_6 + shifted_state16_157_7 + shifted_state16_159_1 + shifted_state16_159_4 + shifted_state16_159_5 + shifted_state16_159_6 + shifted_state16_159_7 + shifted_state16_165_2 + shifted_state16_165_5 + shifted_state16_185_0 + shifted_state16_185_2 + shifted_state16_185_5 + shifted_state16_185_6 + shifted_state16_185_7 + shifted_state16_198_2 + shifted_state16_198_5);
      reservoir_sum_parallel[17] = (shifted_state17_4_1 + shifted_state17_4_2 + shifted_state17_4_5 + shifted_state17_4_6 + shifted_state17_4_7 + shifted_state17_17_1 + shifted_state17_17_2 + shifted_state17_17_4 + shifted_state17_23_0 + shifted_state17_23_2 + shifted_state17_31_0 + shifted_state17_31_1 + shifted_state17_32_2 + shifted_state17_32_3 + shifted_state17_37_0 + shifted_state17_37_1 + shifted_state17_37_2 + shifted_state17_37_3 + shifted_state17_37_4 + shifted_state17_43_5 + shifted_state17_43_6 + shifted_state17_43_7 + shifted_state17_44_3 + shifted_state17_44_4 + shifted_state17_44_5 + shifted_state17_44_6 + shifted_state17_44_7 + shifted_state17_55_0 + shifted_state17_55_1 + shifted_state17_55_5 + shifted_state17_55_6 + shifted_state17_55_7 + shifted_state17_58_3 + shifted_state17_78_0 + shifted_state17_78_2 + shifted_state17_78_3 + shifted_state17_78_4 + shifted_state17_78_6 + shifted_state17_78_7 + shifted_state17_88_0 + shifted_state17_88_2 + shifted_state17_88_3 + shifted_state17_88_4 + shifted_state17_88_7 + shifted_state17_93_0 + shifted_state17_93_3 + shifted_state17_93_4 + shifted_state17_95_2 + shifted_state17_95_4 + shifted_state17_95_6 + shifted_state17_95_7 + shifted_state17_106_1 + shifted_state17_106_3 + shifted_state17_106_4 + shifted_state17_106_5 + shifted_state17_128_0 + shifted_state17_128_3 + shifted_state17_140_1 + shifted_state17_140_2 + shifted_state17_140_3 + shifted_state17_140_4 + shifted_state17_140_5 + shifted_state17_140_7 + shifted_state17_141_0 + shifted_state17_141_1 + shifted_state17_141_2 + shifted_state17_141_3 + shifted_state17_143_1 + shifted_state17_160_0 + shifted_state17_160_1 + shifted_state17_160_2 + shifted_state17_160_5 + shifted_state17_160_6 + shifted_state17_160_7 + shifted_state17_169_0 + shifted_state17_169_1 + shifted_state17_169_4 + shifted_state17_170_1 + shifted_state17_170_3 + shifted_state17_170_4 + shifted_state17_170_5 + shifted_state17_170_6 + shifted_state17_170_7 + shifted_state17_185_3 + shifted_state17_185_5 + shifted_state17_186_0 + shifted_state17_186_4 + shifted_state17_186_5 + shifted_state17_186_6 + shifted_state17_186_7 + shifted_state17_190_1 + shifted_state17_190_3 + shifted_state17_190_5 + shifted_state17_192_0 + shifted_state17_192_1 + shifted_state17_192_2 + shifted_state17_192_5);
      reservoir_sum_parallel[18] = (shifted_state18_3_1 + shifted_state18_3_4 + shifted_state18_3_5 + shifted_state18_3_6 + shifted_state18_3_7 + shifted_state18_4_0 + shifted_state18_4_1 + shifted_state18_4_3 + shifted_state18_4_4 + shifted_state18_4_5 + shifted_state18_4_6 + shifted_state18_4_7 + shifted_state18_7_1 + shifted_state18_7_5 + shifted_state18_7_6 + shifted_state18_7_7 + shifted_state18_10_2 + shifted_state18_22_1 + shifted_state18_27_1 + shifted_state18_27_2 + shifted_state18_27_3 + shifted_state18_27_5 + shifted_state18_27_6 + shifted_state18_27_7 + shifted_state18_47_0 + shifted_state18_47_1 + shifted_state18_47_2 + shifted_state18_67_3 + shifted_state18_67_4 + shifted_state18_78_1 + shifted_state18_82_0 + shifted_state18_82_1 + shifted_state18_82_2 + shifted_state18_82_3 + shifted_state18_82_6 + shifted_state18_86_0 + shifted_state18_86_1 + shifted_state18_86_3 + shifted_state18_86_5 + shifted_state18_86_6 + shifted_state18_86_7 + shifted_state18_100_4 + shifted_state18_113_0 + shifted_state18_113_2 + shifted_state18_113_4 + shifted_state18_113_5 + shifted_state18_113_6 + shifted_state18_113_7 + shifted_state18_116_0 + shifted_state18_116_5 + shifted_state18_121_1 + shifted_state18_121_2 + shifted_state18_121_5 + shifted_state18_123_0 + shifted_state18_123_1 + shifted_state18_123_3 + shifted_state18_123_4 + shifted_state18_123_5 + shifted_state18_123_6 + shifted_state18_123_7 + shifted_state18_135_0 + shifted_state18_135_1 + shifted_state18_135_3 + shifted_state18_135_4 + shifted_state18_135_6 + shifted_state18_135_7 + shifted_state18_139_0 + shifted_state18_139_1 + shifted_state18_139_3 + shifted_state18_143_1 + shifted_state18_143_2 + shifted_state18_143_3 + shifted_state18_143_4 + shifted_state18_151_1 + shifted_state18_151_2 + shifted_state18_151_5 + shifted_state18_151_6 + shifted_state18_151_7 + shifted_state18_153_1 + shifted_state18_153_3 + shifted_state18_153_6 + shifted_state18_153_7 + shifted_state18_164_0 + shifted_state18_164_1 + shifted_state18_164_3 + shifted_state18_166_0 + shifted_state18_166_1 + shifted_state18_166_3 + shifted_state18_166_6 + shifted_state18_166_7 + shifted_state18_173_0 + shifted_state18_173_2 + shifted_state18_173_4 + shifted_state18_173_5 + shifted_state18_173_6 + shifted_state18_173_7 + shifted_state18_180_1 + shifted_state18_180_5 + shifted_state18_180_6 + shifted_state18_180_7 + shifted_state18_188_0 + shifted_state18_188_1 + shifted_state18_188_3 + shifted_state18_188_5 + shifted_state18_188_6 + shifted_state18_188_7 + shifted_state18_196_0 + shifted_state18_196_1 + shifted_state18_196_2 + shifted_state18_196_4 + shifted_state18_196_5 + shifted_state18_196_6 + shifted_state18_196_7);
      reservoir_sum_parallel[19] = (shifted_state19_21_1 + shifted_state19_21_2 + shifted_state19_21_3 + shifted_state19_27_3 + shifted_state19_27_5 + shifted_state19_27_6 + shifted_state19_27_7 + shifted_state19_33_1 + shifted_state19_33_3 + shifted_state19_33_6 + shifted_state19_33_7 + shifted_state19_34_0 + shifted_state19_34_1 + shifted_state19_34_4 + shifted_state19_67_1 + shifted_state19_67_4 + shifted_state19_67_5 + shifted_state19_67_6 + shifted_state19_67_7 + shifted_state19_76_1 + shifted_state19_76_3 + shifted_state19_76_4 + shifted_state19_76_5 + shifted_state19_80_0 + shifted_state19_80_2 + shifted_state19_80_3 + shifted_state19_82_0 + shifted_state19_82_2 + shifted_state19_82_3 + shifted_state19_82_4 + shifted_state19_82_5 + shifted_state19_82_6 + shifted_state19_82_7 + shifted_state19_84_0 + shifted_state19_84_3 + shifted_state19_84_6 + shifted_state19_84_7 + shifted_state19_101_1 + shifted_state19_101_2 + shifted_state19_101_5 + shifted_state19_106_0 + shifted_state19_106_2 + shifted_state19_106_4 + shifted_state19_106_5 + shifted_state19_110_0 + shifted_state19_110_1 + shifted_state19_110_2 + shifted_state19_110_4 + shifted_state19_110_5 + shifted_state19_110_6 + shifted_state19_110_7 + shifted_state19_127_0 + shifted_state19_127_4 + shifted_state19_127_5 + shifted_state19_127_6 + shifted_state19_127_7 + shifted_state19_129_0 + shifted_state19_129_2 + shifted_state19_129_3 + shifted_state19_129_6 + shifted_state19_129_7 + shifted_state19_140_2 + shifted_state19_140_3 + shifted_state19_140_5 + shifted_state19_140_6 + shifted_state19_140_7 + shifted_state19_144_1 + shifted_state19_144_2 + shifted_state19_144_5 + shifted_state19_166_6 + shifted_state19_170_0 + shifted_state19_170_1 + shifted_state19_170_2 + shifted_state19_170_3 + shifted_state19_170_5 + shifted_state19_176_1 + shifted_state19_176_2 + shifted_state19_176_4 + shifted_state19_180_1 + shifted_state19_180_2 + shifted_state19_180_4 + shifted_state19_180_5 + shifted_state19_180_6 + shifted_state19_180_7 + shifted_state19_198_0 + shifted_state19_198_2 + shifted_state19_198_4);
      reservoir_sum_parallel[20] = (shifted_state20_3_2 + shifted_state20_3_3 + shifted_state20_4_0 + shifted_state20_4_1 + shifted_state20_8_1 + shifted_state20_8_3 + shifted_state20_8_4 + shifted_state20_16_1 + shifted_state20_16_3 + shifted_state20_16_4 + shifted_state20_16_5 + shifted_state20_16_6 + shifted_state20_16_7 + shifted_state20_25_3 + shifted_state20_25_5 + shifted_state20_25_6 + shifted_state20_25_7 + shifted_state20_27_0 + shifted_state20_27_2 + shifted_state20_27_4 + shifted_state20_55_1 + shifted_state20_55_4 + shifted_state20_61_1 + shifted_state20_61_3 + shifted_state20_61_6 + shifted_state20_68_4 + shifted_state20_76_0 + shifted_state20_76_4 + shifted_state20_93_0 + shifted_state20_93_1 + shifted_state20_93_2 + shifted_state20_109_2 + shifted_state20_109_4 + shifted_state20_109_5 + shifted_state20_109_6 + shifted_state20_109_7 + shifted_state20_156_1 + shifted_state20_156_2 + shifted_state20_156_3 + shifted_state20_158_0 + shifted_state20_158_3 + shifted_state20_160_1 + shifted_state20_160_2 + shifted_state20_169_0 + shifted_state20_169_2 + shifted_state20_169_3 + shifted_state20_187_1 + shifted_state20_187_3 + shifted_state20_192_0 + shifted_state20_192_3 + shifted_state20_192_4 + shifted_state20_192_6 + shifted_state20_192_7);
      reservoir_sum_parallel[21] = (shifted_state21_7_1 + shifted_state21_7_2 + shifted_state21_7_3 + shifted_state21_7_4 + shifted_state21_7_5 + shifted_state21_7_6 + shifted_state21_7_7 + shifted_state21_22_0 + shifted_state21_22_1 + shifted_state21_22_4 + shifted_state21_26_0 + shifted_state21_26_3 + shifted_state21_27_1 + shifted_state21_27_2 + shifted_state21_27_3 + shifted_state21_27_4 + shifted_state21_27_5 + shifted_state21_27_6 + shifted_state21_27_7 + shifted_state21_32_1 + shifted_state21_32_2 + shifted_state21_32_3 + shifted_state21_32_5 + shifted_state21_32_6 + shifted_state21_32_7 + shifted_state21_34_0 + shifted_state21_34_5 + shifted_state21_34_6 + shifted_state21_34_7 + shifted_state21_37_0 + shifted_state21_37_1 + shifted_state21_37_2 + shifted_state21_37_4 + shifted_state21_55_0 + shifted_state21_55_3 + shifted_state21_75_0 + shifted_state21_75_1 + shifted_state21_75_3 + shifted_state21_75_4 + shifted_state21_100_0 + shifted_state21_100_1 + shifted_state21_100_2 + shifted_state21_100_4 + shifted_state21_100_5 + shifted_state21_100_6 + shifted_state21_100_7 + shifted_state21_109_1 + shifted_state21_109_2 + shifted_state21_109_6 + shifted_state21_109_7 + shifted_state21_113_0 + shifted_state21_113_5 + shifted_state21_113_6 + shifted_state21_113_7 + shifted_state21_116_1 + shifted_state21_116_3 + shifted_state21_116_5 + shifted_state21_116_6 + shifted_state21_116_7 + shifted_state21_124_0 + shifted_state21_124_1 + shifted_state21_124_2 + shifted_state21_124_3 + shifted_state21_124_4 + shifted_state21_124_5 + shifted_state21_124_6 + shifted_state21_124_7 + shifted_state21_134_1 + shifted_state21_134_3 + shifted_state21_134_5 + shifted_state21_134_6 + shifted_state21_134_7 + shifted_state21_140_2 + shifted_state21_140_4 + shifted_state21_140_6 + shifted_state21_140_7 + shifted_state21_150_0 + shifted_state21_150_5 + shifted_state21_150_6 + shifted_state21_150_7 + shifted_state21_158_1 + shifted_state21_158_4 + shifted_state21_158_6 + shifted_state21_158_7 + shifted_state21_162_0 + shifted_state21_162_1 + shifted_state21_162_3 + shifted_state21_166_5 + shifted_state21_172_1 + shifted_state21_172_3 + shifted_state21_172_5 + shifted_state21_172_6 + shifted_state21_172_7 + shifted_state21_177_3 + shifted_state21_177_6 + shifted_state21_177_7 + shifted_state21_180_0 + shifted_state21_180_5);
      reservoir_sum_parallel[22] = (shifted_state22_16_1 + shifted_state22_16_3 + shifted_state22_25_0 + shifted_state22_25_1 + shifted_state22_25_2 + shifted_state22_25_3 + shifted_state22_25_4 + shifted_state22_25_5 + shifted_state22_25_6 + shifted_state22_25_7 + shifted_state22_30_0 + shifted_state22_30_3 + shifted_state22_50_0 + shifted_state22_50_1 + shifted_state22_61_0 + shifted_state22_61_2 + shifted_state22_61_3 + shifted_state22_61_4 + shifted_state22_61_6 + shifted_state22_61_7 + shifted_state22_62_0 + shifted_state22_62_1 + shifted_state22_62_5 + shifted_state22_62_6 + shifted_state22_62_7 + shifted_state22_71_0 + shifted_state22_75_0 + shifted_state22_75_1 + shifted_state22_75_2 + shifted_state22_75_5 + shifted_state22_92_0 + shifted_state22_92_1 + shifted_state22_92_3 + shifted_state22_92_5 + shifted_state22_92_6 + shifted_state22_92_7 + shifted_state22_93_0 + shifted_state22_93_2 + shifted_state22_93_3 + shifted_state22_93_4 + shifted_state22_116_0 + shifted_state22_116_2 + shifted_state22_116_3 + shifted_state22_116_5 + shifted_state22_116_6 + shifted_state22_116_7 + shifted_state22_126_1 + shifted_state22_126_5 + shifted_state22_157_2 + shifted_state22_157_3 + shifted_state22_157_4 + shifted_state22_164_0 + shifted_state22_164_3 + shifted_state22_164_5 + shifted_state22_164_6 + shifted_state22_164_7 + shifted_state22_167_1 + shifted_state22_167_2 + shifted_state22_167_6 + shifted_state22_167_7 + shifted_state22_172_1 + shifted_state22_172_2 + shifted_state22_172_4 + shifted_state22_172_5 + shifted_state22_172_6 + shifted_state22_172_7 + shifted_state22_184_2 + shifted_state22_184_3 + shifted_state22_184_4 + shifted_state22_184_6 + shifted_state22_184_7 + shifted_state22_197_1 + shifted_state22_199_0 + shifted_state22_199_1 + shifted_state22_199_2 + shifted_state22_199_4 + shifted_state22_199_5 + shifted_state22_199_6 + shifted_state22_199_7);
      reservoir_sum_parallel[23] = (shifted_state23_9_0 + shifted_state23_9_1 + shifted_state23_9_2 + shifted_state23_13_2 + shifted_state23_13_4 + shifted_state23_13_5 + shifted_state23_13_6 + shifted_state23_13_7 + shifted_state23_47_0 + shifted_state23_47_3 + shifted_state23_47_5 + shifted_state23_56_0 + shifted_state23_56_3 + shifted_state23_57_2 + shifted_state23_61_2 + shifted_state23_61_5 + shifted_state23_67_0 + shifted_state23_67_1 + shifted_state23_67_4 + shifted_state23_67_5 + shifted_state23_67_6 + shifted_state23_67_7 + shifted_state23_88_2 + shifted_state23_88_5 + shifted_state23_88_6 + shifted_state23_88_7 + shifted_state23_96_0 + shifted_state23_96_1 + shifted_state23_96_3 + shifted_state23_96_4 + shifted_state23_96_5 + shifted_state23_96_6 + shifted_state23_96_7 + shifted_state23_101_2 + shifted_state23_101_3 + shifted_state23_102_1 + shifted_state23_102_4 + shifted_state23_102_6 + shifted_state23_102_7 + shifted_state23_105_0 + shifted_state23_105_3 + shifted_state23_105_4 + shifted_state23_105_6 + shifted_state23_105_7 + shifted_state23_117_2 + shifted_state23_117_4 + shifted_state23_118_4 + shifted_state23_119_1 + shifted_state23_122_0 + shifted_state23_122_1 + shifted_state23_122_3 + shifted_state23_122_5 + shifted_state23_132_1 + shifted_state23_132_2 + shifted_state23_132_3 + shifted_state23_140_0 + shifted_state23_140_2 + shifted_state23_140_5 + shifted_state23_166_1 + shifted_state23_166_2 + shifted_state23_166_5 + shifted_state23_166_6 + shifted_state23_166_7 + shifted_state23_167_1 + shifted_state23_167_3 + shifted_state23_167_4 + shifted_state23_167_5 + shifted_state23_167_6 + shifted_state23_167_7 + shifted_state23_170_2 + shifted_state23_170_3 + shifted_state23_181_0 + shifted_state23_181_2 + shifted_state23_181_3 + shifted_state23_181_4 + shifted_state23_181_5 + shifted_state23_181_6 + shifted_state23_181_7 + shifted_state23_184_0 + shifted_state23_184_1 + shifted_state23_184_4 + shifted_state23_195_2 + shifted_state23_195_3 + shifted_state23_195_4 + shifted_state23_195_6 + shifted_state23_195_7);
      reservoir_sum_parallel[24] = (shifted_state24_1_1 + shifted_state24_1_2 + shifted_state24_1_4 + shifted_state24_1_5 + shifted_state24_1_6 + shifted_state24_1_7 + shifted_state24_3_0 + shifted_state24_3_2 + shifted_state24_3_3 + shifted_state24_3_5 + shifted_state24_3_6 + shifted_state24_3_7 + shifted_state24_9_0 + shifted_state24_9_1 + shifted_state24_9_2 + shifted_state24_9_3 + shifted_state24_9_4 + shifted_state24_9_5 + shifted_state24_9_6 + shifted_state24_9_7 + shifted_state24_13_0 + shifted_state24_13_1 + shifted_state24_13_4 + shifted_state24_13_5 + shifted_state24_13_6 + shifted_state24_13_7 + shifted_state24_22_6 + shifted_state24_22_7 + shifted_state24_29_0 + shifted_state24_29_1 + shifted_state24_29_2 + shifted_state24_32_1 + shifted_state24_32_2 + shifted_state24_32_3 + shifted_state24_32_5 + shifted_state24_32_6 + shifted_state24_32_7 + shifted_state24_38_1 + shifted_state24_38_3 + shifted_state24_49_0 + shifted_state24_49_1 + shifted_state24_49_2 + shifted_state24_49_3 + shifted_state24_49_4 + shifted_state24_63_1 + shifted_state24_63_2 + shifted_state24_69_0 + shifted_state24_69_1 + shifted_state24_69_4 + shifted_state24_69_5 + shifted_state24_69_6 + shifted_state24_69_7 + shifted_state24_87_0 + shifted_state24_87_2 + shifted_state24_87_3 + shifted_state24_87_5 + shifted_state24_87_6 + shifted_state24_87_7 + shifted_state24_96_0 + shifted_state24_96_1 + shifted_state24_96_5 + shifted_state24_96_6 + shifted_state24_96_7 + shifted_state24_102_0 + shifted_state24_102_1 + shifted_state24_102_2 + shifted_state24_102_3 + shifted_state24_102_4 + shifted_state24_102_5 + shifted_state24_102_6 + shifted_state24_102_7 + shifted_state24_116_1 + shifted_state24_116_2 + shifted_state24_116_4 + shifted_state24_131_0 + shifted_state24_131_2 + shifted_state24_131_3 + shifted_state24_131_6 + shifted_state24_131_7 + shifted_state24_154_0 + shifted_state24_154_4 + shifted_state24_154_5 + shifted_state24_154_6 + shifted_state24_154_7 + shifted_state24_169_0 + shifted_state24_169_2 + shifted_state24_169_5 + shifted_state24_169_6 + shifted_state24_169_7 + shifted_state24_178_0 + shifted_state24_180_0 + shifted_state24_180_2 + shifted_state24_180_3 + shifted_state24_180_4 + shifted_state24_180_5 + shifted_state24_180_6 + shifted_state24_180_7);
      reservoir_sum_parallel[25] = (shifted_state25_1_0 + shifted_state25_1_5 + shifted_state25_11_0 + shifted_state25_11_3 + shifted_state25_11_5 + shifted_state25_11_6 + shifted_state25_11_7 + shifted_state25_16_1 + shifted_state25_16_2 + shifted_state25_19_1 + shifted_state25_31_0 + shifted_state25_31_3 + shifted_state25_31_5 + shifted_state25_31_6 + shifted_state25_31_7 + shifted_state25_44_2 + shifted_state25_44_3 + shifted_state25_44_4 + shifted_state25_50_3 + shifted_state25_50_4 + shifted_state25_50_5 + shifted_state25_50_6 + shifted_state25_50_7 + shifted_state25_51_0 + shifted_state25_51_1 + shifted_state25_51_2 + shifted_state25_51_4 + shifted_state25_53_1 + shifted_state25_53_4 + shifted_state25_64_1 + shifted_state25_64_3 + shifted_state25_75_1 + shifted_state25_75_2 + shifted_state25_75_4 + shifted_state25_75_5 + shifted_state25_75_6 + shifted_state25_75_7 + shifted_state25_82_0 + shifted_state25_82_2 + shifted_state25_82_3 + shifted_state25_82_4 + shifted_state25_82_5 + shifted_state25_82_6 + shifted_state25_82_7 + shifted_state25_83_1 + shifted_state25_83_4 + shifted_state25_98_4 + shifted_state25_109_0 + shifted_state25_109_1 + shifted_state25_109_2 + shifted_state25_122_1 + shifted_state25_122_2 + shifted_state25_122_4 + shifted_state25_145_0 + shifted_state25_145_4 + shifted_state25_153_0 + shifted_state25_153_2 + shifted_state25_153_4 + shifted_state25_153_5 + shifted_state25_153_6 + shifted_state25_153_7 + shifted_state25_157_2 + shifted_state25_157_3 + shifted_state25_162_0 + shifted_state25_162_2 + shifted_state25_170_3 + shifted_state25_170_5 + shifted_state25_185_0 + shifted_state25_185_1 + shifted_state25_185_4 + shifted_state25_187_0 + shifted_state25_187_2 + shifted_state25_187_4 + shifted_state25_187_5 + shifted_state25_187_6 + shifted_state25_187_7 + shifted_state25_192_1 + shifted_state25_192_3 + shifted_state25_195_0 + shifted_state25_195_1 + shifted_state25_195_3);
      reservoir_sum_parallel[26] = (shifted_state26_3_0 + shifted_state26_3_2 + shifted_state26_3_3 + shifted_state26_3_4 + shifted_state26_11_2 + shifted_state26_11_4 + shifted_state26_18_0 + shifted_state26_18_1 + shifted_state26_18_3 + shifted_state26_27_0 + shifted_state26_27_2 + shifted_state26_27_4 + shifted_state26_27_5 + shifted_state26_27_6 + shifted_state26_27_7 + shifted_state26_30_0 + shifted_state26_30_1 + shifted_state26_30_4 + shifted_state26_30_6 + shifted_state26_30_7 + shifted_state26_33_0 + shifted_state26_33_2 + shifted_state26_33_3 + shifted_state26_36_2 + shifted_state26_36_3 + shifted_state26_54_4 + shifted_state26_54_6 + shifted_state26_58_0 + shifted_state26_58_1 + shifted_state26_58_3 + shifted_state26_58_5 + shifted_state26_58_6 + shifted_state26_58_7 + shifted_state26_89_0 + shifted_state26_89_2 + shifted_state26_89_3 + shifted_state26_89_5 + shifted_state26_89_6 + shifted_state26_89_7 + shifted_state26_100_0 + shifted_state26_100_3 + shifted_state26_117_0 + shifted_state26_117_1 + shifted_state26_117_2 + shifted_state26_117_4 + shifted_state26_117_6 + shifted_state26_117_7 + shifted_state26_168_0 + shifted_state26_168_2 + shifted_state26_168_3 + shifted_state26_168_5 + shifted_state26_168_6 + shifted_state26_168_7 + shifted_state26_185_3 + shifted_state26_185_4 + shifted_state26_185_5 + shifted_state26_185_6 + shifted_state26_185_7);
      reservoir_sum_parallel[27] = (shifted_state27_2_0 + shifted_state27_2_4 + shifted_state27_22_0 + shifted_state27_22_1 + shifted_state27_22_2 + shifted_state27_22_4 + shifted_state27_22_5 + shifted_state27_22_6 + shifted_state27_22_7 + shifted_state27_24_1 + shifted_state27_24_2 + shifted_state27_24_4 + shifted_state27_25_0 + shifted_state27_25_2 + shifted_state27_25_4 + shifted_state27_27_1 + shifted_state27_27_2 + shifted_state27_46_1 + shifted_state27_65_1 + shifted_state27_65_2 + shifted_state27_65_3 + shifted_state27_65_5 + shifted_state27_65_6 + shifted_state27_65_7 + shifted_state27_89_1 + shifted_state27_89_4 + shifted_state27_104_0 + shifted_state27_104_5 + shifted_state27_104_6 + shifted_state27_104_7 + shifted_state27_107_0 + shifted_state27_107_1 + shifted_state27_107_2 + shifted_state27_109_0 + shifted_state27_109_1 + shifted_state27_114_3 + shifted_state27_114_4 + shifted_state27_114_5 + shifted_state27_114_6 + shifted_state27_114_7 + shifted_state27_117_1 + shifted_state27_117_4 + shifted_state27_117_5 + shifted_state27_117_6 + shifted_state27_117_7 + shifted_state27_127_2 + shifted_state27_127_4 + shifted_state27_127_6 + shifted_state27_127_7 + shifted_state27_132_0 + shifted_state27_132_1 + shifted_state27_132_3 + shifted_state27_132_4 + shifted_state27_132_5 + shifted_state27_140_2 + shifted_state27_140_4 + shifted_state27_140_5 + shifted_state27_140_7 + shifted_state27_148_4 + shifted_state27_148_5 + shifted_state27_148_6 + shifted_state27_148_7 + shifted_state27_155_1 + shifted_state27_155_2 + shifted_state27_155_3 + shifted_state27_155_4 + shifted_state27_167_0 + shifted_state27_175_1 + shifted_state27_175_3 + shifted_state27_175_5 + shifted_state27_175_6 + shifted_state27_175_7 + shifted_state27_176_3 + shifted_state27_176_4 + shifted_state27_176_5 + shifted_state27_176_6 + shifted_state27_176_7 + shifted_state27_184_1 + shifted_state27_184_2 + shifted_state27_191_1 + shifted_state27_191_4 + shifted_state27_191_5 + shifted_state27_191_6 + shifted_state27_191_7 + shifted_state27_193_0 + shifted_state27_193_1 + shifted_state27_193_4);
      reservoir_sum_parallel[28] = (shifted_state28_1_0 + shifted_state28_1_1 + shifted_state28_1_2 + shifted_state28_1_4 + shifted_state28_1_6 + shifted_state28_1_7 + shifted_state28_2_0 + shifted_state28_2_1 + shifted_state28_2_4 + shifted_state28_2_5 + shifted_state28_2_6 + shifted_state28_2_7 + shifted_state28_4_2 + shifted_state28_4_3 + shifted_state28_9_5 + shifted_state28_9_6 + shifted_state28_9_7 + shifted_state28_24_0 + shifted_state28_24_1 + shifted_state28_24_3 + shifted_state28_24_4 + shifted_state28_42_0 + shifted_state28_42_1 + shifted_state28_42_3 + shifted_state28_42_4 + shifted_state28_42_5 + shifted_state28_42_6 + shifted_state28_42_7 + shifted_state28_46_0 + shifted_state28_46_1 + shifted_state28_46_2 + shifted_state28_46_3 + shifted_state28_46_4 + shifted_state28_46_5 + shifted_state28_46_6 + shifted_state28_46_7 + shifted_state28_71_3 + shifted_state28_71_4 + shifted_state28_72_2 + shifted_state28_72_3 + shifted_state28_72_4 + shifted_state28_72_5 + shifted_state28_72_7 + shifted_state28_76_1 + shifted_state28_76_2 + shifted_state28_76_3 + shifted_state28_76_4 + shifted_state28_76_5 + shifted_state28_76_6 + shifted_state28_76_7 + shifted_state28_79_0 + shifted_state28_79_1 + shifted_state28_80_2 + shifted_state28_80_3 + shifted_state28_97_0 + shifted_state28_97_2 + shifted_state28_97_3 + shifted_state28_97_4 + shifted_state28_100_0 + shifted_state28_100_1 + shifted_state28_100_2 + shifted_state28_100_5 + shifted_state28_100_6 + shifted_state28_100_7 + shifted_state28_105_0 + shifted_state28_105_3 + shifted_state28_105_4 + shifted_state28_105_5 + shifted_state28_107_0 + shifted_state28_107_2 + shifted_state28_107_4 + shifted_state28_107_5 + shifted_state28_121_0 + shifted_state28_121_5 + shifted_state28_136_0 + shifted_state28_136_1 + shifted_state28_136_4 + shifted_state28_136_5 + shifted_state28_136_6 + shifted_state28_136_7 + shifted_state28_140_0 + shifted_state28_140_2 + shifted_state28_140_4 + shifted_state28_140_5 + shifted_state28_140_6 + shifted_state28_140_7 + shifted_state28_141_3 + shifted_state28_141_4 + shifted_state28_144_1 + shifted_state28_144_3 + shifted_state28_144_6 + shifted_state28_144_7 + shifted_state28_170_1 + shifted_state28_170_2 + shifted_state28_170_3 + shifted_state28_170_4 + shifted_state28_172_0 + shifted_state28_172_4 + shifted_state28_186_0 + shifted_state28_186_2 + shifted_state28_186_4 + shifted_state28_186_5 + shifted_state28_186_6 + shifted_state28_186_7 + shifted_state28_187_0 + shifted_state28_187_1 + shifted_state28_187_2 + shifted_state28_187_6 + shifted_state28_187_7 + shifted_state28_189_4 + shifted_state28_189_6 + shifted_state28_189_7 + shifted_state28_195_2 + shifted_state28_195_4 + shifted_state28_198_0 + shifted_state28_198_4 + shifted_state28_198_5 + shifted_state28_198_6 + shifted_state28_198_7);
      reservoir_sum_parallel[29] = (shifted_state29_0_0 + shifted_state29_0_2 + shifted_state29_0_3 + shifted_state29_0_4 + shifted_state29_0_6 + shifted_state29_0_7 + shifted_state29_14_1 + shifted_state29_14_2 + shifted_state29_14_3 + shifted_state29_14_5 + shifted_state29_14_6 + shifted_state29_14_7 + shifted_state29_16_0 + shifted_state29_16_2 + shifted_state29_16_4 + shifted_state29_16_5 + shifted_state29_16_6 + shifted_state29_16_7 + shifted_state29_18_3 + shifted_state29_18_5 + shifted_state29_18_6 + shifted_state29_18_7 + shifted_state29_28_1 + shifted_state29_28_5 + shifted_state29_35_2 + shifted_state29_35_3 + shifted_state29_35_5 + shifted_state29_35_6 + shifted_state29_35_7 + shifted_state29_49_1 + shifted_state29_49_2 + shifted_state29_49_5 + shifted_state29_49_6 + shifted_state29_49_7 + shifted_state29_60_0 + shifted_state29_60_2 + shifted_state29_60_4 + shifted_state29_63_1 + shifted_state29_63_2 + shifted_state29_63_4 + shifted_state29_63_5 + shifted_state29_63_6 + shifted_state29_63_7 + shifted_state29_78_0 + shifted_state29_78_1 + shifted_state29_78_3 + shifted_state29_78_4 + shifted_state29_78_5 + shifted_state29_78_6 + shifted_state29_78_7 + shifted_state29_96_3 + shifted_state29_96_5 + shifted_state29_96_6 + shifted_state29_96_7 + shifted_state29_106_0 + shifted_state29_106_1 + shifted_state29_106_3 + shifted_state29_107_3 + shifted_state29_107_5 + shifted_state29_107_6 + shifted_state29_107_7 + shifted_state29_127_0 + shifted_state29_127_1 + shifted_state29_127_4 + shifted_state29_127_6 + shifted_state29_127_7 + shifted_state29_171_0 + shifted_state29_171_1 + shifted_state29_171_2 + shifted_state29_171_4 + shifted_state29_171_5 + shifted_state29_171_6 + shifted_state29_171_7 + shifted_state29_177_3 + shifted_state29_177_5 + shifted_state29_177_6 + shifted_state29_177_7 + shifted_state29_183_0 + shifted_state29_183_2 + shifted_state29_183_3 + shifted_state29_183_4 + shifted_state29_183_5 + shifted_state29_183_6 + shifted_state29_183_7 + shifted_state29_190_0 + shifted_state29_190_2 + shifted_state29_190_3 + shifted_state29_191_0 + shifted_state29_191_1 + shifted_state29_191_4 + shifted_state29_191_5 + shifted_state29_191_6 + shifted_state29_191_7 + shifted_state29_196_1 + shifted_state29_196_4 + shifted_state29_199_3 + shifted_state29_199_5 + shifted_state29_199_6 + shifted_state29_199_7);
      reservoir_sum_parallel[30] = (shifted_state30_7_3 + shifted_state30_8_2 + shifted_state30_8_3 + shifted_state30_18_0 + shifted_state30_18_2 + shifted_state30_18_4 + shifted_state30_18_5 + shifted_state30_18_6 + shifted_state30_18_7 + shifted_state30_53_0 + shifted_state30_53_2 + shifted_state30_53_4 + shifted_state30_53_6 + shifted_state30_53_7 + shifted_state30_62_0 + shifted_state30_62_2 + shifted_state30_62_3 + shifted_state30_62_4 + shifted_state30_62_6 + shifted_state30_62_7 + shifted_state30_64_5 + shifted_state30_71_0 + shifted_state30_71_1 + shifted_state30_71_2 + shifted_state30_71_3 + shifted_state30_77_0 + shifted_state30_77_1 + shifted_state30_77_2 + shifted_state30_77_4 + shifted_state30_91_4 + shifted_state30_104_0 + shifted_state30_104_1 + shifted_state30_104_2 + shifted_state30_104_4 + shifted_state30_104_5 + shifted_state30_104_6 + shifted_state30_104_7 + shifted_state30_107_1 + shifted_state30_107_5 + shifted_state30_107_6 + shifted_state30_107_7 + shifted_state30_115_0 + shifted_state30_115_2 + shifted_state30_117_0 + shifted_state30_117_1 + shifted_state30_117_4 + shifted_state30_117_5 + shifted_state30_117_6 + shifted_state30_117_7 + shifted_state30_120_3 + shifted_state30_120_4 + shifted_state30_120_5 + shifted_state30_120_6 + shifted_state30_120_7 + shifted_state30_129_0 + shifted_state30_129_3 + shifted_state30_142_0 + shifted_state30_142_1 + shifted_state30_142_2 + shifted_state30_142_3 + shifted_state30_142_5 + shifted_state30_142_6 + shifted_state30_142_7 + shifted_state30_151_0 + shifted_state30_151_1 + shifted_state30_151_3 + shifted_state30_151_4 + shifted_state30_151_5 + shifted_state30_151_6 + shifted_state30_151_7 + shifted_state30_156_0 + shifted_state30_156_2 + shifted_state30_156_3 + shifted_state30_156_4 + shifted_state30_156_6 + shifted_state30_156_7 + shifted_state30_162_0 + shifted_state30_162_4 + shifted_state30_162_5 + shifted_state30_169_0 + shifted_state30_169_2 + shifted_state30_169_3 + shifted_state30_169_4 + shifted_state30_169_6 + shifted_state30_169_7 + shifted_state30_184_0 + shifted_state30_184_3 + shifted_state30_186_0 + shifted_state30_186_3 + shifted_state30_186_4 + shifted_state30_186_5 + shifted_state30_186_6 + shifted_state30_186_7 + shifted_state30_188_0 + shifted_state30_188_2 + shifted_state30_188_3 + shifted_state30_188_4);
      reservoir_sum_parallel[31] = (shifted_state31_11_0 + shifted_state31_11_2 + shifted_state31_25_1 + shifted_state31_25_3 + shifted_state31_52_0 + shifted_state31_52_2 + shifted_state31_52_3 + shifted_state31_52_6 + shifted_state31_56_0 + shifted_state31_56_1 + shifted_state31_56_3 + shifted_state31_56_4 + shifted_state31_56_6 + shifted_state31_56_7 + shifted_state31_58_0 + shifted_state31_58_1 + shifted_state31_58_2 + shifted_state31_58_3 + shifted_state31_58_5 + shifted_state31_58_6 + shifted_state31_58_7 + shifted_state31_61_0 + shifted_state31_61_1 + shifted_state31_61_2 + shifted_state31_61_6 + shifted_state31_62_0 + shifted_state31_62_5 + shifted_state31_101_0 + shifted_state31_101_5 + shifted_state31_106_0 + shifted_state31_106_1 + shifted_state31_106_2 + shifted_state31_106_4 + shifted_state31_111_1 + shifted_state31_111_2 + shifted_state31_111_5 + shifted_state31_111_6 + shifted_state31_111_7 + shifted_state31_120_0 + shifted_state31_120_2 + shifted_state31_129_0 + shifted_state31_129_2 + shifted_state31_129_5 + shifted_state31_129_6 + shifted_state31_129_7 + shifted_state31_139_1 + shifted_state31_139_4 + shifted_state31_139_5 + shifted_state31_139_6 + shifted_state31_139_7 + shifted_state31_145_2 + shifted_state31_145_5 + shifted_state31_145_6 + shifted_state31_145_7 + shifted_state31_149_0 + shifted_state31_149_1 + shifted_state31_149_3 + shifted_state31_155_0 + shifted_state31_155_3 + shifted_state31_155_4 + shifted_state31_155_5 + shifted_state31_174_5 + shifted_state31_174_6 + shifted_state31_174_7 + shifted_state31_178_2 + shifted_state31_178_4 + shifted_state31_178_5 + shifted_state31_178_6 + shifted_state31_178_7 + shifted_state31_179_0 + shifted_state31_179_1 + shifted_state31_179_2 + shifted_state31_179_3 + shifted_state31_179_4 + shifted_state31_179_5 + shifted_state31_179_6 + shifted_state31_179_7 + shifted_state31_182_0 + shifted_state31_182_2 + shifted_state31_182_3 + shifted_state31_182_4 + shifted_state31_182_5 + shifted_state31_182_6 + shifted_state31_182_7 + shifted_state31_194_0 + shifted_state31_194_2 + shifted_state31_194_3 + shifted_state31_194_5 + shifted_state31_194_6 + shifted_state31_194_7);
      reservoir_sum_parallel[32] = (shifted_state32_3_3 + shifted_state32_4_1 + shifted_state32_4_3 + shifted_state32_4_5 + shifted_state32_4_6 + shifted_state32_4_7 + shifted_state32_9_1 + shifted_state32_9_4 + shifted_state32_14_0 + shifted_state32_14_2 + shifted_state32_22_0 + shifted_state32_22_2 + shifted_state32_39_0 + shifted_state32_39_1 + shifted_state32_39_2 + shifted_state32_39_3 + shifted_state32_39_4 + shifted_state32_39_5 + shifted_state32_39_6 + shifted_state32_39_7 + shifted_state32_46_1 + shifted_state32_46_2 + shifted_state32_46_4 + shifted_state32_46_5 + shifted_state32_46_6 + shifted_state32_46_7 + shifted_state32_57_0 + shifted_state32_57_4 + shifted_state32_61_2 + shifted_state32_61_6 + shifted_state32_72_4 + shifted_state32_72_5 + shifted_state32_72_6 + shifted_state32_72_7 + shifted_state32_102_0 + shifted_state32_102_3 + shifted_state32_109_0 + shifted_state32_109_2 + shifted_state32_109_3 + shifted_state32_109_5 + shifted_state32_124_0 + shifted_state32_124_3 + shifted_state32_124_4 + shifted_state32_124_6 + shifted_state32_124_7 + shifted_state32_126_0 + shifted_state32_126_1 + shifted_state32_126_3 + shifted_state32_126_4 + shifted_state32_126_6 + shifted_state32_126_7 + shifted_state32_133_0 + shifted_state32_133_1 + shifted_state32_133_2 + shifted_state32_133_3 + shifted_state32_133_4 + shifted_state32_133_5 + shifted_state32_133_6 + shifted_state32_133_7 + shifted_state32_138_0 + shifted_state32_138_4 + shifted_state32_138_6 + shifted_state32_138_7 + shifted_state32_161_0 + shifted_state32_161_1 + shifted_state32_161_5 + shifted_state32_161_6 + shifted_state32_161_7 + shifted_state32_172_1 + shifted_state32_172_6 + shifted_state32_191_1 + shifted_state32_191_4 + shifted_state32_191_5 + shifted_state32_198_0 + shifted_state32_198_1 + shifted_state32_198_3 + shifted_state32_198_4 + shifted_state32_198_5);
      reservoir_sum_parallel[33] = (shifted_state33_2_0 + shifted_state33_2_1 + shifted_state33_2_2 + shifted_state33_2_3 + shifted_state33_8_0 + shifted_state33_8_3 + shifted_state33_9_1 + shifted_state33_9_3 + shifted_state33_9_4 + shifted_state33_9_5 + shifted_state33_9_6 + shifted_state33_9_7 + shifted_state33_17_0 + shifted_state33_17_2 + shifted_state33_17_3 + shifted_state33_17_4 + shifted_state33_17_5 + shifted_state33_17_6 + shifted_state33_17_7 + shifted_state33_34_1 + shifted_state33_34_2 + shifted_state33_38_0 + shifted_state33_38_3 + shifted_state33_38_4 + shifted_state33_38_5 + shifted_state33_38_6 + shifted_state33_38_7 + shifted_state33_51_0 + shifted_state33_51_2 + shifted_state33_51_5 + shifted_state33_51_6 + shifted_state33_51_7 + shifted_state33_57_0 + shifted_state33_57_4 + shifted_state33_59_0 + shifted_state33_59_3 + shifted_state33_59_4 + shifted_state33_79_0 + shifted_state33_79_2 + shifted_state33_79_3 + shifted_state33_79_4 + shifted_state33_79_5 + shifted_state33_79_6 + shifted_state33_79_7 + shifted_state33_106_1 + shifted_state33_108_1 + shifted_state33_108_2 + shifted_state33_108_3 + shifted_state33_108_5 + shifted_state33_108_6 + shifted_state33_108_7 + shifted_state33_129_0 + shifted_state33_129_1 + shifted_state33_129_4 + shifted_state33_131_1 + shifted_state33_131_3 + shifted_state33_131_5 + shifted_state33_141_1 + shifted_state33_141_3 + shifted_state33_141_4 + shifted_state33_141_6 + shifted_state33_141_7 + shifted_state33_155_1 + shifted_state33_155_2 + shifted_state33_155_3 + shifted_state33_155_5 + shifted_state33_155_6 + shifted_state33_155_7 + shifted_state33_164_5 + shifted_state33_168_0 + shifted_state33_168_5 + shifted_state33_168_6 + shifted_state33_168_7 + shifted_state33_173_1 + shifted_state33_173_2 + shifted_state33_173_3 + shifted_state33_173_4 + shifted_state33_173_5 + shifted_state33_173_6 + shifted_state33_173_7 + shifted_state33_177_3 + shifted_state33_178_0 + shifted_state33_178_1 + shifted_state33_178_3 + shifted_state33_178_4 + shifted_state33_178_5 + shifted_state33_178_6 + shifted_state33_178_7 + shifted_state33_179_1 + shifted_state33_179_3 + shifted_state33_179_5 + shifted_state33_184_0 + shifted_state33_184_4 + shifted_state33_184_5);
      reservoir_sum_parallel[34] = (shifted_state34_5_0 + shifted_state34_5_1 + shifted_state34_34_1 + shifted_state34_34_3 + shifted_state34_34_6 + shifted_state34_34_7 + shifted_state34_36_0 + shifted_state34_36_2 + shifted_state34_36_4 + shifted_state34_36_5 + shifted_state34_36_6 + shifted_state34_36_7 + shifted_state34_41_0 + shifted_state34_41_1 + shifted_state34_41_2 + shifted_state34_41_3 + shifted_state34_41_4 + shifted_state34_41_5 + shifted_state34_41_7 + shifted_state34_46_0 + shifted_state34_46_2 + shifted_state34_46_3 + shifted_state34_46_4 + shifted_state34_63_2 + shifted_state34_63_5 + shifted_state34_80_0 + shifted_state34_80_2 + shifted_state34_80_4 + shifted_state34_90_1 + shifted_state34_90_2 + shifted_state34_90_5 + shifted_state34_92_2 + shifted_state34_92_5 + shifted_state34_99_1 + shifted_state34_99_2 + shifted_state34_99_3 + shifted_state34_99_4 + shifted_state34_99_5 + shifted_state34_99_6 + shifted_state34_99_7 + shifted_state34_101_0 + shifted_state34_106_0 + shifted_state34_106_3 + shifted_state34_106_5 + shifted_state34_107_0 + shifted_state34_107_2 + shifted_state34_107_4 + shifted_state34_108_3 + shifted_state34_108_4 + shifted_state34_108_5 + shifted_state34_120_1 + shifted_state34_120_2 + shifted_state34_120_3 + shifted_state34_120_4 + shifted_state34_138_0 + shifted_state34_138_1 + shifted_state34_138_2 + shifted_state34_138_5 + shifted_state34_138_6 + shifted_state34_138_7 + shifted_state34_148_0 + shifted_state34_148_2 + shifted_state34_148_3 + shifted_state34_148_5 + shifted_state34_148_6 + shifted_state34_148_7 + shifted_state34_152_0 + shifted_state34_152_1 + shifted_state34_162_0 + shifted_state34_162_1 + shifted_state34_162_2 + shifted_state34_163_1 + shifted_state34_163_2 + shifted_state34_163_4 + shifted_state34_163_5 + shifted_state34_163_6 + shifted_state34_163_7 + shifted_state34_186_1 + shifted_state34_186_4 + shifted_state34_186_5 + shifted_state34_186_6 + shifted_state34_186_7 + shifted_state34_195_1 + shifted_state34_195_4);
      reservoir_sum_parallel[35] = (shifted_state35_2_1 + shifted_state35_2_2 + shifted_state35_2_4 + shifted_state35_23_0 + shifted_state35_23_1 + shifted_state35_23_5 + shifted_state35_30_1 + shifted_state35_30_2 + shifted_state35_37_0 + shifted_state35_42_0 + shifted_state35_42_1 + shifted_state35_42_3 + shifted_state35_56_0 + shifted_state35_56_1 + shifted_state35_56_5 + shifted_state35_56_6 + shifted_state35_56_7 + shifted_state35_59_0 + shifted_state35_59_2 + shifted_state35_64_0 + shifted_state35_64_4 + shifted_state35_64_6 + shifted_state35_64_7 + shifted_state35_81_0 + shifted_state35_81_1 + shifted_state35_81_4 + shifted_state35_88_2 + shifted_state35_96_0 + shifted_state35_96_1 + shifted_state35_96_2 + shifted_state35_96_5 + shifted_state35_100_0 + shifted_state35_100_3 + shifted_state35_100_4 + shifted_state35_100_6 + shifted_state35_100_7 + shifted_state35_102_0 + shifted_state35_102_1 + shifted_state35_102_2 + shifted_state35_102_5 + shifted_state35_102_6 + shifted_state35_102_7 + shifted_state35_105_1 + shifted_state35_105_2 + shifted_state35_122_2 + shifted_state35_122_3 + shifted_state35_122_5 + shifted_state35_122_6 + shifted_state35_122_7 + shifted_state35_133_0 + shifted_state35_133_1 + shifted_state35_133_5 + shifted_state35_133_6 + shifted_state35_133_7 + shifted_state35_142_1 + shifted_state35_145_0 + shifted_state35_145_3 + shifted_state35_157_0 + shifted_state35_157_1 + shifted_state35_157_2 + shifted_state35_157_4 + shifted_state35_157_6 + shifted_state35_157_7 + shifted_state35_165_1 + shifted_state35_165_3 + shifted_state35_165_4 + shifted_state35_165_5 + shifted_state35_165_6 + shifted_state35_165_7 + shifted_state35_173_3 + shifted_state35_173_4 + shifted_state35_173_5 + shifted_state35_174_0 + shifted_state35_174_1 + shifted_state35_174_3 + shifted_state35_174_6 + shifted_state35_174_7 + shifted_state35_183_2 + shifted_state35_186_0 + shifted_state35_186_1 + shifted_state35_186_3 + shifted_state35_186_4 + shifted_state35_186_5 + shifted_state35_186_6 + shifted_state35_186_7 + shifted_state35_187_1 + shifted_state35_187_3 + shifted_state35_187_5 + shifted_state35_187_6 + shifted_state35_187_7 + shifted_state35_191_0 + shifted_state35_191_2 + shifted_state35_191_4 + shifted_state35_191_5);
      reservoir_sum_parallel[36] = (shifted_state36_0_2 + shifted_state36_0_4 + shifted_state36_16_0 + shifted_state36_16_1 + shifted_state36_32_0 + shifted_state36_32_1 + shifted_state36_32_3 + shifted_state36_32_4 + shifted_state36_32_5 + shifted_state36_32_6 + shifted_state36_32_7 + shifted_state36_35_3 + shifted_state36_35_4 + shifted_state36_39_1 + shifted_state36_39_2 + shifted_state36_39_3 + shifted_state36_39_4 + shifted_state36_39_5 + shifted_state36_39_6 + shifted_state36_39_7 + shifted_state36_44_1 + shifted_state36_44_2 + shifted_state36_44_4 + shifted_state36_50_0 + shifted_state36_50_3 + shifted_state36_50_4 + shifted_state36_55_1 + shifted_state36_55_5 + shifted_state36_55_6 + shifted_state36_55_7 + shifted_state36_70_1 + shifted_state36_70_4 + shifted_state36_70_5 + shifted_state36_76_0 + shifted_state36_76_1 + shifted_state36_76_4 + shifted_state36_76_5 + shifted_state36_76_6 + shifted_state36_76_7 + shifted_state36_97_0 + shifted_state36_97_3 + shifted_state36_97_4 + shifted_state36_97_5 + shifted_state36_97_6 + shifted_state36_97_7 + shifted_state36_105_0 + shifted_state36_105_3 + shifted_state36_105_4 + shifted_state36_105_5 + shifted_state36_134_1 + shifted_state36_137_0 + shifted_state36_137_3 + shifted_state36_137_4 + shifted_state36_137_5 + shifted_state36_137_6 + shifted_state36_137_7 + shifted_state36_143_0 + shifted_state36_143_3 + shifted_state36_143_4 + shifted_state36_155_2 + shifted_state36_155_4 + shifted_state36_155_5 + shifted_state36_155_6 + shifted_state36_155_7 + shifted_state36_160_0 + shifted_state36_160_3 + shifted_state36_160_4 + shifted_state36_160_5 + shifted_state36_160_6 + shifted_state36_160_7 + shifted_state36_163_0 + shifted_state36_163_1 + shifted_state36_163_2 + shifted_state36_163_3 + shifted_state36_193_0 + shifted_state36_193_2 + shifted_state36_193_4 + shifted_state36_193_6 + shifted_state36_193_7);
      reservoir_sum_parallel[37] = (shifted_state37_4_0 + shifted_state37_33_1 + shifted_state37_33_3 + shifted_state37_33_4 + shifted_state37_33_5 + shifted_state37_33_6 + shifted_state37_33_7 + shifted_state37_38_1 + shifted_state37_38_3 + shifted_state37_38_4 + shifted_state37_38_6 + shifted_state37_38_7 + shifted_state37_66_5 + shifted_state37_81_0 + shifted_state37_81_4 + shifted_state37_88_0 + shifted_state37_88_1 + shifted_state37_88_4 + shifted_state37_88_6 + shifted_state37_88_7 + shifted_state37_89_0 + shifted_state37_89_1 + shifted_state37_89_2 + shifted_state37_89_3 + shifted_state37_89_4 + shifted_state37_89_6 + shifted_state37_89_7 + shifted_state37_98_0 + shifted_state37_98_2 + shifted_state37_98_4 + shifted_state37_121_0 + shifted_state37_121_1 + shifted_state37_121_3 + shifted_state37_150_1 + shifted_state37_150_3 + shifted_state37_150_4 + shifted_state37_158_0 + shifted_state37_158_2 + shifted_state37_165_1 + shifted_state37_165_2 + shifted_state37_165_3 + shifted_state37_165_4 + shifted_state37_165_5 + shifted_state37_165_6 + shifted_state37_165_7 + shifted_state37_173_0 + shifted_state37_173_2 + shifted_state37_173_3 + shifted_state37_173_4 + shifted_state37_173_5 + shifted_state37_173_6 + shifted_state37_173_7 + shifted_state37_185_4 + shifted_state37_185_6 + shifted_state37_185_7 + shifted_state37_186_0 + shifted_state37_186_1 + shifted_state37_186_3 + shifted_state37_186_4 + shifted_state37_186_5 + shifted_state37_186_6 + shifted_state37_186_7 + shifted_state37_187_1 + shifted_state37_187_3 + shifted_state37_187_4 + shifted_state37_187_5 + shifted_state37_187_6 + shifted_state37_187_7 + shifted_state37_191_5 + shifted_state37_191_6 + shifted_state37_191_7);
      reservoir_sum_parallel[38] = (shifted_state38_9_0 + shifted_state38_9_3 + shifted_state38_9_4 + shifted_state38_9_6 + shifted_state38_9_7 + shifted_state38_13_0 + shifted_state38_13_1 + shifted_state38_13_2 + shifted_state38_13_4 + shifted_state38_13_6 + shifted_state38_13_7 + shifted_state38_41_0 + shifted_state38_41_1 + shifted_state38_41_4 + shifted_state38_41_5 + shifted_state38_41_6 + shifted_state38_41_7 + shifted_state38_42_1 + shifted_state38_42_2 + shifted_state38_42_4 + shifted_state38_45_0 + shifted_state38_45_1 + shifted_state38_45_2 + shifted_state38_45_3 + shifted_state38_45_4 + shifted_state38_45_6 + shifted_state38_45_7 + shifted_state38_72_0 + shifted_state38_72_1 + shifted_state38_72_3 + shifted_state38_72_4 + shifted_state38_72_5 + shifted_state38_72_6 + shifted_state38_72_7 + shifted_state38_76_2 + shifted_state38_76_3 + shifted_state38_76_4 + shifted_state38_76_5 + shifted_state38_76_6 + shifted_state38_76_7 + shifted_state38_83_0 + shifted_state38_83_1 + shifted_state38_83_2 + shifted_state38_87_4 + shifted_state38_87_5 + shifted_state38_87_6 + shifted_state38_87_7 + shifted_state38_103_0 + shifted_state38_103_1 + shifted_state38_103_2 + shifted_state38_103_4 + shifted_state38_120_0 + shifted_state38_120_2 + shifted_state38_120_3 + shifted_state38_124_0 + shifted_state38_124_2 + shifted_state38_124_4 + shifted_state38_124_5 + shifted_state38_135_0 + shifted_state38_135_1 + shifted_state38_135_3 + shifted_state38_135_5 + shifted_state38_157_0 + shifted_state38_157_1 + shifted_state38_157_3 + shifted_state38_162_1 + shifted_state38_162_3 + shifted_state38_162_4 + shifted_state38_162_5 + shifted_state38_162_6 + shifted_state38_162_7 + shifted_state38_167_1 + shifted_state38_167_3 + shifted_state38_167_4 + shifted_state38_172_0 + shifted_state38_172_1 + shifted_state38_172_3 + shifted_state38_172_4 + shifted_state38_172_5 + shifted_state38_172_6 + shifted_state38_172_7 + shifted_state38_175_2 + shifted_state38_179_1 + shifted_state38_179_2 + shifted_state38_179_3);
      reservoir_sum_parallel[39] = (shifted_state39_1_0 + shifted_state39_1_2 + shifted_state39_1_3 + shifted_state39_1_4 + shifted_state39_1_6 + shifted_state39_1_7 + shifted_state39_3_0 + shifted_state39_3_2 + shifted_state39_3_3 + shifted_state39_3_5 + shifted_state39_20_3 + shifted_state39_20_5 + shifted_state39_26_1 + shifted_state39_26_4 + shifted_state39_34_0 + shifted_state39_34_2 + shifted_state39_43_0 + shifted_state39_43_3 + shifted_state39_43_6 + shifted_state39_69_1 + shifted_state39_69_2 + shifted_state39_69_4 + shifted_state39_69_5 + shifted_state39_69_6 + shifted_state39_69_7 + shifted_state39_80_0 + shifted_state39_80_1 + shifted_state39_80_3 + shifted_state39_85_0 + shifted_state39_85_2 + shifted_state39_85_4 + shifted_state39_85_5 + shifted_state39_85_6 + shifted_state39_85_7 + shifted_state39_86_3 + shifted_state39_86_4 + shifted_state39_86_5 + shifted_state39_86_6 + shifted_state39_86_7 + shifted_state39_88_0 + shifted_state39_88_1 + shifted_state39_88_2 + shifted_state39_88_4 + shifted_state39_95_1 + shifted_state39_95_3 + shifted_state39_95_4 + shifted_state39_95_5 + shifted_state39_95_6 + shifted_state39_95_7 + shifted_state39_105_0 + shifted_state39_105_2 + shifted_state39_105_3 + shifted_state39_105_4 + shifted_state39_105_5 + shifted_state39_105_6 + shifted_state39_105_7 + shifted_state39_106_0 + shifted_state39_106_1 + shifted_state39_106_2 + shifted_state39_106_3 + shifted_state39_106_4 + shifted_state39_106_5 + shifted_state39_106_6 + shifted_state39_106_7 + shifted_state39_115_0 + shifted_state39_115_1 + shifted_state39_115_2 + shifted_state39_121_2 + shifted_state39_121_3 + shifted_state39_121_5 + shifted_state39_121_6 + shifted_state39_121_7 + shifted_state39_132_4 + shifted_state39_161_1 + shifted_state39_161_2 + shifted_state39_161_5 + shifted_state39_161_6 + shifted_state39_161_7 + shifted_state39_162_0 + shifted_state39_162_2 + shifted_state39_162_3 + shifted_state39_162_4 + shifted_state39_169_0 + shifted_state39_169_3 + shifted_state39_169_5 + shifted_state39_172_0 + shifted_state39_172_1 + shifted_state39_172_2 + shifted_state39_172_4 + shifted_state39_172_6 + shifted_state39_172_7 + shifted_state39_175_0 + shifted_state39_175_1 + shifted_state39_175_2 + shifted_state39_175_3 + shifted_state39_175_4 + shifted_state39_175_5 + shifted_state39_175_6 + shifted_state39_175_7 + shifted_state39_176_1 + shifted_state39_176_2 + shifted_state39_176_4 + shifted_state39_176_6 + shifted_state39_176_7 + shifted_state39_187_1);
      reservoir_sum_parallel[40] = (shifted_state40_6_0 + shifted_state40_6_1 + shifted_state40_6_5 + shifted_state40_6_6 + shifted_state40_6_7 + shifted_state40_9_0 + shifted_state40_9_2 + shifted_state40_9_3 + shifted_state40_9_5 + shifted_state40_9_6 + shifted_state40_9_7 + shifted_state40_21_1 + shifted_state40_21_3 + shifted_state40_21_4 + shifted_state40_21_5 + shifted_state40_21_6 + shifted_state40_21_7 + shifted_state40_23_0 + shifted_state40_23_3 + shifted_state40_23_5 + shifted_state40_23_6 + shifted_state40_23_7 + shifted_state40_35_5 + shifted_state40_41_0 + shifted_state40_41_2 + shifted_state40_41_3 + shifted_state40_41_4 + shifted_state40_41_5 + shifted_state40_41_6 + shifted_state40_41_7 + shifted_state40_46_0 + shifted_state40_48_1 + shifted_state40_48_4 + shifted_state40_48_5 + shifted_state40_49_0 + shifted_state40_57_0 + shifted_state40_57_3 + shifted_state40_57_4 + shifted_state40_75_3 + shifted_state40_75_4 + shifted_state40_75_5 + shifted_state40_75_6 + shifted_state40_75_7 + shifted_state40_77_0 + shifted_state40_77_1 + shifted_state40_77_2 + shifted_state40_89_0 + shifted_state40_89_1 + shifted_state40_89_2 + shifted_state40_89_3 + shifted_state40_89_4 + shifted_state40_89_5 + shifted_state40_89_6 + shifted_state40_89_7 + shifted_state40_112_0 + shifted_state40_112_4 + shifted_state40_112_5 + shifted_state40_112_6 + shifted_state40_112_7 + shifted_state40_119_5 + shifted_state40_119_6 + shifted_state40_119_7 + shifted_state40_120_0 + shifted_state40_120_1 + shifted_state40_120_3 + shifted_state40_120_5 + shifted_state40_120_6 + shifted_state40_120_7 + shifted_state40_123_0 + shifted_state40_123_1 + shifted_state40_123_2 + shifted_state40_123_3 + shifted_state40_123_4 + shifted_state40_123_5 + shifted_state40_123_6 + shifted_state40_123_7 + shifted_state40_126_0 + shifted_state40_126_1 + shifted_state40_126_2 + shifted_state40_126_4 + shifted_state40_126_5 + shifted_state40_126_6 + shifted_state40_126_7 + shifted_state40_138_3 + shifted_state40_138_4 + shifted_state40_138_5 + shifted_state40_138_6 + shifted_state40_138_7 + shifted_state40_153_0 + shifted_state40_153_1 + shifted_state40_153_2 + shifted_state40_153_5 + shifted_state40_153_6 + shifted_state40_153_7 + shifted_state40_156_0 + shifted_state40_156_2 + shifted_state40_156_3 + shifted_state40_156_4 + shifted_state40_156_5 + shifted_state40_156_6 + shifted_state40_156_7 + shifted_state40_177_0 + shifted_state40_177_1 + shifted_state40_177_3 + shifted_state40_177_4);
      reservoir_sum_parallel[41] = (shifted_state41_31_2 + shifted_state41_31_4 + shifted_state41_31_5 + shifted_state41_31_6 + shifted_state41_31_7 + shifted_state41_43_0 + shifted_state41_43_2 + shifted_state41_43_3 + shifted_state41_43_4 + shifted_state41_43_5 + shifted_state41_43_6 + shifted_state41_43_7 + shifted_state41_50_0 + shifted_state41_50_1 + shifted_state41_50_2 + shifted_state41_50_3 + shifted_state41_50_5 + shifted_state41_50_6 + shifted_state41_50_7 + shifted_state41_53_0 + shifted_state41_53_2 + shifted_state41_53_3 + shifted_state41_53_4 + shifted_state41_53_6 + shifted_state41_53_7 + shifted_state41_74_1 + shifted_state41_74_2 + shifted_state41_74_4 + shifted_state41_83_0 + shifted_state41_83_1 + shifted_state41_83_3 + shifted_state41_83_5 + shifted_state41_83_6 + shifted_state41_83_7 + shifted_state41_97_0 + shifted_state41_97_1 + shifted_state41_97_5 + shifted_state41_97_6 + shifted_state41_97_7 + shifted_state41_103_0 + shifted_state41_103_1 + shifted_state41_104_0 + shifted_state41_104_1 + shifted_state41_104_2 + shifted_state41_104_4 + shifted_state41_112_2 + shifted_state41_112_4 + shifted_state41_112_5 + shifted_state41_124_0 + shifted_state41_124_1 + shifted_state41_124_4 + shifted_state41_147_4 + shifted_state41_147_5 + shifted_state41_167_1 + shifted_state41_167_2 + shifted_state41_167_3 + shifted_state41_167_4 + shifted_state41_168_0 + shifted_state41_168_3 + shifted_state41_168_4 + shifted_state41_168_5 + shifted_state41_168_6 + shifted_state41_168_7 + shifted_state41_173_0 + shifted_state41_173_1 + shifted_state41_173_3 + shifted_state41_173_4 + shifted_state41_173_5 + shifted_state41_173_7 + shifted_state41_179_0 + shifted_state41_179_2 + shifted_state41_179_3 + shifted_state41_179_4 + shifted_state41_179_5 + shifted_state41_179_6 + shifted_state41_179_7 + shifted_state41_195_3 + shifted_state41_195_4 + shifted_state41_195_6 + shifted_state41_195_7);
      reservoir_sum_parallel[42] = (shifted_state42_26_0 + shifted_state42_26_1 + shifted_state42_26_4 + shifted_state42_26_5 + shifted_state42_26_6 + shifted_state42_26_7 + shifted_state42_42_1 + shifted_state42_42_2 + shifted_state42_42_3 + shifted_state42_42_5 + shifted_state42_43_0 + shifted_state42_43_3 + shifted_state42_43_5 + shifted_state42_43_6 + shifted_state42_43_7 + shifted_state42_74_2 + shifted_state42_74_6 + shifted_state42_74_7 + shifted_state42_82_1 + shifted_state42_82_2 + shifted_state42_82_4 + shifted_state42_85_0 + shifted_state42_85_5 + shifted_state42_95_1 + shifted_state42_95_2 + shifted_state42_95_3 + shifted_state42_95_4 + shifted_state42_95_5 + shifted_state42_95_6 + shifted_state42_95_7 + shifted_state42_139_0 + shifted_state42_139_1 + shifted_state42_139_2 + shifted_state42_139_3 + shifted_state42_143_0 + shifted_state42_143_1 + shifted_state42_143_4 + shifted_state42_143_6 + shifted_state42_143_7 + shifted_state42_153_1 + shifted_state42_153_3 + shifted_state42_153_4 + shifted_state42_167_5 + shifted_state42_198_0 + shifted_state42_198_1 + shifted_state42_198_2 + shifted_state42_198_3 + shifted_state42_198_4);
      reservoir_sum_parallel[43] = (shifted_state43_7_1 + shifted_state43_7_3 + shifted_state43_7_4 + shifted_state43_7_5 + shifted_state43_7_6 + shifted_state43_7_7 + shifted_state43_22_0 + shifted_state43_22_1 + shifted_state43_22_3 + shifted_state43_22_5 + shifted_state43_55_1 + shifted_state43_55_5 + shifted_state43_93_0 + shifted_state43_93_3 + shifted_state43_93_4 + shifted_state43_106_1 + shifted_state43_106_5 + shifted_state43_106_6 + shifted_state43_106_7 + shifted_state43_109_1 + shifted_state43_109_3 + shifted_state43_109_5 + shifted_state43_109_6 + shifted_state43_109_7 + shifted_state43_130_1 + shifted_state43_130_3 + shifted_state43_135_1 + shifted_state43_135_2 + shifted_state43_135_4 + shifted_state43_135_5 + shifted_state43_135_6 + shifted_state43_135_7 + shifted_state43_158_0 + shifted_state43_158_1 + shifted_state43_158_2 + shifted_state43_158_4 + shifted_state43_173_1 + shifted_state43_173_2 + shifted_state43_173_4 + shifted_state43_185_1 + shifted_state43_185_5 + shifted_state43_185_6 + shifted_state43_185_7);
      reservoir_sum_parallel[44] = (shifted_state44_3_0 + shifted_state44_3_1 + shifted_state44_3_3 + shifted_state44_3_5 + shifted_state44_3_6 + shifted_state44_3_7 + shifted_state44_16_0 + shifted_state44_16_3 + shifted_state44_16_4 + shifted_state44_16_6 + shifted_state44_16_7 + shifted_state44_20_0 + shifted_state44_20_1 + shifted_state44_20_3 + shifted_state44_55_0 + shifted_state44_55_1 + shifted_state44_55_3 + shifted_state44_55_4 + shifted_state44_63_0 + shifted_state44_63_1 + shifted_state44_63_2 + shifted_state44_63_3 + shifted_state44_63_6 + shifted_state44_63_7 + shifted_state44_68_0 + shifted_state44_68_1 + shifted_state44_68_3 + shifted_state44_68_4 + shifted_state44_68_5 + shifted_state44_68_6 + shifted_state44_68_7 + shifted_state44_69_0 + shifted_state44_69_1 + shifted_state44_69_4 + shifted_state44_69_5 + shifted_state44_69_6 + shifted_state44_69_7 + shifted_state44_70_1 + shifted_state44_71_1 + shifted_state44_71_2 + shifted_state44_71_4 + shifted_state44_72_1 + shifted_state44_72_3 + shifted_state44_72_5 + shifted_state44_79_2 + shifted_state44_79_4 + shifted_state44_79_5 + shifted_state44_79_6 + shifted_state44_79_7 + shifted_state44_81_3 + shifted_state44_87_2 + shifted_state44_87_3 + shifted_state44_87_5 + shifted_state44_87_6 + shifted_state44_87_7 + shifted_state44_91_1 + shifted_state44_91_4 + shifted_state44_108_1 + shifted_state44_108_2 + shifted_state44_129_2 + shifted_state44_129_5 + shifted_state44_136_0 + shifted_state44_136_1 + shifted_state44_136_5 + shifted_state44_136_6 + shifted_state44_136_7 + shifted_state44_147_5 + shifted_state44_150_2 + shifted_state44_172_0 + shifted_state44_172_4 + shifted_state44_174_1 + shifted_state44_174_2 + shifted_state44_174_3 + shifted_state44_174_5 + shifted_state44_174_6 + shifted_state44_174_7 + shifted_state44_186_2 + shifted_state44_186_4 + shifted_state44_186_5 + shifted_state44_186_6 + shifted_state44_186_7 + shifted_state44_193_0 + shifted_state44_193_2 + shifted_state44_193_5 + shifted_state44_193_6 + shifted_state44_193_7);
      reservoir_sum_parallel[45] = (shifted_state45_29_0 + shifted_state45_29_1 + shifted_state45_29_2 + shifted_state45_29_3 + shifted_state45_33_1 + shifted_state45_33_2 + shifted_state45_33_3 + shifted_state45_44_1 + shifted_state45_44_3 + shifted_state45_44_6 + shifted_state45_54_1 + shifted_state45_54_2 + shifted_state45_54_3 + shifted_state45_54_5 + shifted_state45_55_0 + shifted_state45_55_1 + shifted_state45_55_2 + shifted_state45_55_3 + shifted_state45_55_4 + shifted_state45_55_6 + shifted_state45_55_7 + shifted_state45_58_0 + shifted_state45_58_2 + shifted_state45_58_3 + shifted_state45_58_5 + shifted_state45_58_6 + shifted_state45_58_7 + shifted_state45_71_1 + shifted_state45_71_2 + shifted_state45_71_5 + shifted_state45_71_6 + shifted_state45_71_7 + shifted_state45_74_2 + shifted_state45_74_4 + shifted_state45_78_0 + shifted_state45_78_2 + shifted_state45_78_3 + shifted_state45_79_0 + shifted_state45_79_1 + shifted_state45_79_2 + shifted_state45_79_4 + shifted_state45_82_0 + shifted_state45_82_2 + shifted_state45_82_3 + shifted_state45_82_4 + shifted_state45_82_6 + shifted_state45_82_7 + shifted_state45_85_4 + shifted_state45_86_0 + shifted_state45_86_2 + shifted_state45_86_3 + shifted_state45_86_4 + shifted_state45_86_5 + shifted_state45_86_6 + shifted_state45_86_7 + shifted_state45_91_0 + shifted_state45_91_2 + shifted_state45_91_3 + shifted_state45_91_4 + shifted_state45_91_6 + shifted_state45_91_7 + shifted_state45_99_0 + shifted_state45_99_2 + shifted_state45_99_3 + shifted_state45_99_5 + shifted_state45_121_0 + shifted_state45_121_1 + shifted_state45_121_2 + shifted_state45_121_4 + shifted_state45_121_5 + shifted_state45_121_6 + shifted_state45_121_7 + shifted_state45_124_0 + shifted_state45_124_1 + shifted_state45_124_2 + shifted_state45_124_4 + shifted_state45_124_5 + shifted_state45_132_0 + shifted_state45_132_2 + shifted_state45_132_3 + shifted_state45_133_3 + shifted_state45_133_4 + shifted_state45_133_5 + shifted_state45_157_4 + shifted_state45_164_0 + shifted_state45_164_3 + shifted_state45_164_5 + shifted_state45_174_0 + shifted_state45_174_2 + shifted_state45_174_3 + shifted_state45_174_5 + shifted_state45_174_6 + shifted_state45_174_7 + shifted_state45_192_0 + shifted_state45_192_1 + shifted_state45_192_3 + shifted_state45_192_4 + shifted_state45_195_1 + shifted_state45_195_3 + shifted_state45_195_5 + shifted_state45_195_6 + shifted_state45_195_7 + shifted_state45_197_1 + shifted_state45_197_3 + shifted_state45_197_5 + shifted_state45_197_6 + shifted_state45_197_7);
      reservoir_sum_parallel[46] = (shifted_state46_33_5 + shifted_state46_40_0 + shifted_state46_40_2 + shifted_state46_40_4 + shifted_state46_42_1 + shifted_state46_42_2 + shifted_state46_42_5 + shifted_state46_59_1 + shifted_state46_59_2 + shifted_state46_59_5 + shifted_state46_59_6 + shifted_state46_59_7 + shifted_state46_61_0 + shifted_state46_61_5 + shifted_state46_68_3 + shifted_state46_68_6 + shifted_state46_68_7 + shifted_state46_91_4 + shifted_state46_91_5 + shifted_state46_91_6 + shifted_state46_91_7 + shifted_state46_93_1 + shifted_state46_93_3 + shifted_state46_93_5 + shifted_state46_93_6 + shifted_state46_93_7 + shifted_state46_106_0 + shifted_state46_106_1 + shifted_state46_106_4 + shifted_state46_106_5 + shifted_state46_106_6 + shifted_state46_106_7 + shifted_state46_109_0 + shifted_state46_109_1 + shifted_state46_109_2 + shifted_state46_109_3 + shifted_state46_116_1 + shifted_state46_116_3 + shifted_state46_123_2 + shifted_state46_123_3 + shifted_state46_123_4 + shifted_state46_123_5 + shifted_state46_123_6 + shifted_state46_123_7 + shifted_state46_125_1 + shifted_state46_126_0 + shifted_state46_126_4 + shifted_state46_126_5 + shifted_state46_126_6 + shifted_state46_126_7 + shifted_state46_136_3 + shifted_state46_136_4 + shifted_state46_136_5 + shifted_state46_136_6 + shifted_state46_136_7 + shifted_state46_138_0 + shifted_state46_138_1 + shifted_state46_138_2 + shifted_state46_138_3 + shifted_state46_138_5 + shifted_state46_146_0 + shifted_state46_146_1 + shifted_state46_146_3 + shifted_state46_146_5 + shifted_state46_146_6 + shifted_state46_146_7 + shifted_state46_147_1 + shifted_state46_147_2 + shifted_state46_147_6 + shifted_state46_149_0 + shifted_state46_149_3 + shifted_state46_149_6 + shifted_state46_149_7 + shifted_state46_174_0 + shifted_state46_174_2 + shifted_state46_174_4 + shifted_state46_181_2 + shifted_state46_181_4 + shifted_state46_184_1 + shifted_state46_184_2 + shifted_state46_184_4 + shifted_state46_184_5 + shifted_state46_184_6 + shifted_state46_184_7);
      reservoir_sum_parallel[47] = (shifted_state47_11_0 + shifted_state47_11_3 + shifted_state47_11_4 + shifted_state47_19_0 + shifted_state47_19_2 + shifted_state47_19_3 + shifted_state47_32_1 + shifted_state47_32_2 + shifted_state47_32_3 + shifted_state47_32_4 + shifted_state47_32_5 + shifted_state47_32_6 + shifted_state47_32_7 + shifted_state47_53_3 + shifted_state47_53_4 + shifted_state47_53_5 + shifted_state47_63_0 + shifted_state47_63_2 + shifted_state47_63_3 + shifted_state47_63_4 + shifted_state47_63_5 + shifted_state47_63_6 + shifted_state47_63_7 + shifted_state47_72_1 + shifted_state47_72_3 + shifted_state47_72_4 + shifted_state47_72_5 + shifted_state47_72_6 + shifted_state47_72_7 + shifted_state47_73_0 + shifted_state47_73_1 + shifted_state47_73_2 + shifted_state47_73_6 + shifted_state47_73_7 + shifted_state47_85_5 + shifted_state47_93_1 + shifted_state47_93_3 + shifted_state47_93_5 + shifted_state47_93_6 + shifted_state47_93_7 + shifted_state47_98_0 + shifted_state47_98_1 + shifted_state47_98_2 + shifted_state47_98_3 + shifted_state47_98_4 + shifted_state47_98_5 + shifted_state47_98_6 + shifted_state47_98_7 + shifted_state47_100_1 + shifted_state47_100_3 + shifted_state47_105_1 + shifted_state47_105_4 + shifted_state47_105_5 + shifted_state47_105_6 + shifted_state47_105_7 + shifted_state47_137_1 + shifted_state47_137_5 + shifted_state47_137_6 + shifted_state47_137_7 + shifted_state47_146_1 + shifted_state47_146_2 + shifted_state47_146_4 + shifted_state47_146_5 + shifted_state47_146_6 + shifted_state47_146_7 + shifted_state47_150_0 + shifted_state47_150_5 + shifted_state47_150_6 + shifted_state47_150_7 + shifted_state47_159_0 + shifted_state47_159_5 + shifted_state47_185_2 + shifted_state47_185_5 + shifted_state47_185_6 + shifted_state47_185_7 + shifted_state47_188_3 + shifted_state47_188_4 + shifted_state47_188_5 + shifted_state47_188_6 + shifted_state47_188_7 + shifted_state47_199_1);
      reservoir_sum_parallel[48] = (shifted_state48_8_2 + shifted_state48_8_4 + shifted_state48_8_5 + shifted_state48_8_6 + shifted_state48_8_7 + shifted_state48_25_0 + shifted_state48_25_2 + shifted_state48_32_0 + shifted_state48_32_4 + shifted_state48_32_5 + shifted_state48_32_6 + shifted_state48_32_7 + shifted_state48_35_1 + shifted_state48_35_4 + shifted_state48_35_5 + shifted_state48_38_1 + shifted_state48_38_2 + shifted_state48_61_1 + shifted_state48_61_2 + shifted_state48_61_4 + shifted_state48_61_5 + shifted_state48_62_0 + shifted_state48_62_1 + shifted_state48_62_2 + shifted_state48_62_3 + shifted_state48_62_4 + shifted_state48_62_6 + shifted_state48_62_7 + shifted_state48_70_1 + shifted_state48_70_3 + shifted_state48_70_6 + shifted_state48_70_7 + shifted_state48_77_1 + shifted_state48_77_5 + shifted_state48_78_2 + shifted_state48_78_4 + shifted_state48_78_5 + shifted_state48_78_6 + shifted_state48_78_7 + shifted_state48_94_0 + shifted_state48_94_1 + shifted_state48_94_2 + shifted_state48_94_3 + shifted_state48_94_4 + shifted_state48_94_5 + shifted_state48_94_6 + shifted_state48_94_7 + shifted_state48_102_1 + shifted_state48_102_5 + shifted_state48_117_1 + shifted_state48_117_2 + shifted_state48_117_3 + shifted_state48_125_0 + shifted_state48_125_2 + shifted_state48_125_3 + shifted_state48_133_0 + shifted_state48_133_3 + shifted_state48_133_5 + shifted_state48_141_0 + shifted_state48_141_2 + shifted_state48_141_3 + shifted_state48_141_4 + shifted_state48_141_6 + shifted_state48_141_7 + shifted_state48_148_0 + shifted_state48_148_2 + shifted_state48_148_3 + shifted_state48_155_0 + shifted_state48_155_1 + shifted_state48_155_3 + shifted_state48_155_4 + shifted_state48_155_5 + shifted_state48_155_6 + shifted_state48_155_7 + shifted_state48_163_3 + shifted_state48_163_5 + shifted_state48_163_6 + shifted_state48_163_7 + shifted_state48_173_0 + shifted_state48_173_2 + shifted_state48_173_5 + shifted_state48_173_6 + shifted_state48_173_7 + shifted_state48_178_1 + shifted_state48_178_2 + shifted_state48_178_4 + shifted_state48_178_5 + shifted_state48_178_6 + shifted_state48_178_7 + shifted_state48_187_0 + shifted_state48_187_1 + shifted_state48_187_2 + shifted_state48_187_3 + shifted_state48_187_4 + shifted_state48_187_5 + shifted_state48_187_6 + shifted_state48_187_7 + shifted_state48_190_0 + shifted_state48_190_1 + shifted_state48_190_3 + shifted_state48_190_4);
      reservoir_sum_parallel[49] = (shifted_state49_4_0 + shifted_state49_4_1 + shifted_state49_4_2 + shifted_state49_4_3 + shifted_state49_4_4 + shifted_state49_4_6 + shifted_state49_4_7 + shifted_state49_34_3 + shifted_state49_34_4 + shifted_state49_34_5 + shifted_state49_34_6 + shifted_state49_34_7 + shifted_state49_38_0 + shifted_state49_38_3 + shifted_state49_53_0 + shifted_state49_53_2 + shifted_state49_62_1 + shifted_state49_62_3 + shifted_state49_62_4 + shifted_state49_74_1 + shifted_state49_74_2 + shifted_state49_74_3 + shifted_state49_74_4 + shifted_state49_74_5 + shifted_state49_74_6 + shifted_state49_74_7 + shifted_state49_99_1 + shifted_state49_99_2 + shifted_state49_99_3 + shifted_state49_109_1 + shifted_state49_109_3 + shifted_state49_109_5 + shifted_state49_132_3 + shifted_state49_132_4 + shifted_state49_132_6 + shifted_state49_132_7 + shifted_state49_145_0 + shifted_state49_145_2 + shifted_state49_145_4 + shifted_state49_157_1 + shifted_state49_157_3 + shifted_state49_157_5 + shifted_state49_157_6 + shifted_state49_157_7 + shifted_state49_159_0 + shifted_state49_159_1 + shifted_state49_159_2);
      reservoir_sum_parallel[50] = (shifted_state50_23_2 + shifted_state50_23_3 + shifted_state50_59_2 + shifted_state50_59_4 + shifted_state50_59_5 + shifted_state50_59_6 + shifted_state50_59_7 + shifted_state50_61_0 + shifted_state50_61_1 + shifted_state50_61_2 + shifted_state50_61_5 + shifted_state50_61_6 + shifted_state50_61_7 + shifted_state50_66_1 + shifted_state50_66_2 + shifted_state50_66_3 + shifted_state50_66_5 + shifted_state50_77_0 + shifted_state50_77_2 + shifted_state50_77_3 + shifted_state50_77_5 + shifted_state50_77_6 + shifted_state50_77_7 + shifted_state50_81_1 + shifted_state50_81_4 + shifted_state50_83_0 + shifted_state50_83_3 + shifted_state50_83_5 + shifted_state50_95_1 + shifted_state50_95_2 + shifted_state50_95_3 + shifted_state50_95_4 + shifted_state50_95_5 + shifted_state50_95_6 + shifted_state50_95_7 + shifted_state50_100_0 + shifted_state50_100_2 + shifted_state50_100_3 + shifted_state50_100_4 + shifted_state50_100_6 + shifted_state50_100_7 + shifted_state50_110_1 + shifted_state50_110_2 + shifted_state50_110_5 + shifted_state50_110_6 + shifted_state50_110_7 + shifted_state50_114_3 + shifted_state50_139_2 + shifted_state50_139_5 + shifted_state50_139_6 + shifted_state50_139_7 + shifted_state50_150_1 + shifted_state50_150_2 + shifted_state50_150_3 + shifted_state50_161_2 + shifted_state50_161_3 + shifted_state50_161_6 + shifted_state50_161_7 + shifted_state50_164_0 + shifted_state50_164_3 + shifted_state50_164_5 + shifted_state50_164_6 + shifted_state50_164_7 + shifted_state50_169_1 + shifted_state50_169_4 + shifted_state50_169_5 + shifted_state50_169_6 + shifted_state50_169_7 + shifted_state50_170_0 + shifted_state50_170_4 + shifted_state50_178_1 + shifted_state50_178_2 + shifted_state50_178_3 + shifted_state50_178_5 + shifted_state50_178_6 + shifted_state50_178_7);
      reservoir_sum_parallel[51] = (shifted_state51_19_0 + shifted_state51_19_2 + shifted_state51_19_3 + shifted_state51_20_0 + shifted_state51_20_5 + shifted_state51_20_6 + shifted_state51_20_7 + shifted_state51_58_2 + shifted_state51_58_5 + shifted_state51_59_0 + shifted_state51_59_1 + shifted_state51_59_2 + shifted_state51_59_4 + shifted_state51_66_0 + shifted_state51_66_2 + shifted_state51_66_3 + shifted_state51_66_5 + shifted_state51_66_6 + shifted_state51_66_7 + shifted_state51_99_0 + shifted_state51_99_3 + shifted_state51_99_4 + shifted_state51_99_5 + shifted_state51_99_6 + shifted_state51_99_7 + shifted_state51_108_2 + shifted_state51_108_3 + shifted_state51_108_4 + shifted_state51_108_5 + shifted_state51_108_6 + shifted_state51_108_7 + shifted_state51_157_2 + shifted_state51_190_0 + shifted_state51_190_1 + shifted_state51_190_2 + shifted_state51_190_3 + shifted_state51_198_1 + shifted_state51_198_2 + shifted_state51_198_3 + shifted_state51_198_4 + shifted_state51_198_5 + shifted_state51_198_6 + shifted_state51_198_7 + shifted_state51_199_1 + shifted_state51_199_2 + shifted_state51_199_4);
      reservoir_sum_parallel[52] = (shifted_state52_9_0 + shifted_state52_9_1 + shifted_state52_9_2 + shifted_state52_9_4 + shifted_state52_9_5 + shifted_state52_9_6 + shifted_state52_9_7 + shifted_state52_26_3 + shifted_state52_26_5 + shifted_state52_26_6 + shifted_state52_26_7 + shifted_state52_48_1 + shifted_state52_48_2 + shifted_state52_48_3 + shifted_state52_48_5 + shifted_state52_53_5 + shifted_state52_53_6 + shifted_state52_53_7 + shifted_state52_71_0 + shifted_state52_71_3 + shifted_state52_71_5 + shifted_state52_71_6 + shifted_state52_71_7 + shifted_state52_79_0 + shifted_state52_79_1 + shifted_state52_79_3 + shifted_state52_79_4 + shifted_state52_79_5 + shifted_state52_79_6 + shifted_state52_79_7 + shifted_state52_86_0 + shifted_state52_86_1 + shifted_state52_86_3 + shifted_state52_86_6 + shifted_state52_86_7 + shifted_state52_94_1 + shifted_state52_94_3 + shifted_state52_94_4 + shifted_state52_112_1 + shifted_state52_112_3 + shifted_state52_119_0 + shifted_state52_119_2 + shifted_state52_119_5 + shifted_state52_119_6 + shifted_state52_119_7 + shifted_state52_142_0 + shifted_state52_142_1 + shifted_state52_142_2 + shifted_state52_142_5 + shifted_state52_144_0 + shifted_state52_144_3 + shifted_state52_144_5 + shifted_state52_151_1 + shifted_state52_151_2 + shifted_state52_151_3 + shifted_state52_151_5 + shifted_state52_174_3 + shifted_state52_174_4 + shifted_state52_174_5 + shifted_state52_174_6 + shifted_state52_174_7 + shifted_state52_180_2 + shifted_state52_180_3 + shifted_state52_180_4 + shifted_state52_180_5 + shifted_state52_180_6 + shifted_state52_180_7 + shifted_state52_184_0 + shifted_state52_184_2 + shifted_state52_184_3 + shifted_state52_184_4 + shifted_state52_189_1 + shifted_state52_189_3 + shifted_state52_199_1 + shifted_state52_199_2);
      reservoir_sum_parallel[53] = (shifted_state53_1_3 + shifted_state53_6_0 + shifted_state53_6_2 + shifted_state53_11_0 + shifted_state53_11_4 + shifted_state53_11_6 + shifted_state53_11_7 + shifted_state53_13_2 + shifted_state53_13_4 + shifted_state53_13_6 + shifted_state53_13_7 + shifted_state53_20_1 + shifted_state53_20_2 + shifted_state53_20_4 + shifted_state53_24_2 + shifted_state53_24_3 + shifted_state53_24_5 + shifted_state53_24_6 + shifted_state53_24_7 + shifted_state53_25_0 + shifted_state53_25_3 + shifted_state53_25_4 + shifted_state53_25_6 + shifted_state53_25_7 + shifted_state53_27_1 + shifted_state53_27_2 + shifted_state53_27_3 + shifted_state53_27_4 + shifted_state53_27_5 + shifted_state53_29_1 + shifted_state53_29_2 + shifted_state53_29_3 + shifted_state53_29_4 + shifted_state53_29_6 + shifted_state53_29_7 + shifted_state53_30_0 + shifted_state53_30_2 + shifted_state53_30_3 + shifted_state53_30_4 + shifted_state53_30_5 + shifted_state53_30_6 + shifted_state53_30_7 + shifted_state53_37_0 + shifted_state53_37_1 + shifted_state53_37_2 + shifted_state53_51_0 + shifted_state53_51_1 + shifted_state53_64_1 + shifted_state53_64_3 + shifted_state53_64_5 + shifted_state53_64_6 + shifted_state53_64_7 + shifted_state53_74_1 + shifted_state53_74_2 + shifted_state53_74_6 + shifted_state53_74_7 + shifted_state53_140_2 + shifted_state53_140_4 + shifted_state53_140_5 + shifted_state53_141_1 + shifted_state53_141_2 + shifted_state53_141_3 + shifted_state53_142_2 + shifted_state53_142_3 + shifted_state53_142_4 + shifted_state53_142_5 + shifted_state53_142_7 + shifted_state53_148_2 + shifted_state53_148_3 + shifted_state53_148_5 + shifted_state53_148_6 + shifted_state53_148_7 + shifted_state53_154_4 + shifted_state53_167_0 + shifted_state53_167_1 + shifted_state53_167_2 + shifted_state53_167_3 + shifted_state53_167_4 + shifted_state53_167_5 + shifted_state53_167_7 + shifted_state53_189_0 + shifted_state53_189_1 + shifted_state53_189_2 + shifted_state53_189_3 + shifted_state53_189_5 + shifted_state53_191_1 + shifted_state53_191_2 + shifted_state53_191_3 + shifted_state53_191_4 + shifted_state53_191_5 + shifted_state53_191_6 + shifted_state53_191_7);
      reservoir_sum_parallel[54] = (shifted_state54_23_1 + shifted_state54_23_4 + shifted_state54_23_5 + shifted_state54_23_6 + shifted_state54_23_7 + shifted_state54_24_1 + shifted_state54_24_3 + shifted_state54_24_4 + shifted_state54_24_5 + shifted_state54_24_6 + shifted_state54_24_7 + shifted_state54_28_0 + shifted_state54_28_3 + shifted_state54_31_0 + shifted_state54_31_5 + shifted_state54_38_0 + shifted_state54_38_1 + shifted_state54_38_3 + shifted_state54_38_4 + shifted_state54_55_5 + shifted_state54_55_6 + shifted_state54_55_7 + shifted_state54_56_1 + shifted_state54_56_2 + shifted_state54_56_3 + shifted_state54_59_1 + shifted_state54_59_4 + shifted_state54_59_6 + shifted_state54_59_7 + shifted_state54_70_2 + shifted_state54_70_3 + shifted_state54_82_0 + shifted_state54_82_2 + shifted_state54_82_4 + shifted_state54_82_5 + shifted_state54_96_0 + shifted_state54_96_2 + shifted_state54_96_4 + shifted_state54_96_6 + shifted_state54_96_7 + shifted_state54_110_1 + shifted_state54_110_4 + shifted_state54_110_5 + shifted_state54_110_6 + shifted_state54_110_7 + shifted_state54_115_0 + shifted_state54_115_1 + shifted_state54_115_2 + shifted_state54_115_3 + shifted_state54_130_0 + shifted_state54_136_0 + shifted_state54_136_3 + shifted_state54_140_1 + shifted_state54_140_2 + shifted_state54_140_4 + shifted_state54_156_1 + shifted_state54_156_2 + shifted_state54_156_4 + shifted_state54_156_5 + shifted_state54_156_6 + shifted_state54_156_7 + shifted_state54_161_1 + shifted_state54_161_4 + shifted_state54_161_5 + shifted_state54_161_6 + shifted_state54_161_7 + shifted_state54_188_0 + shifted_state54_188_2 + shifted_state54_188_3 + shifted_state54_189_2 + shifted_state54_189_3 + shifted_state54_193_2 + shifted_state54_193_4 + shifted_state54_193_5 + shifted_state54_195_0 + shifted_state54_195_1 + shifted_state54_195_2 + shifted_state54_195_3 + shifted_state54_195_4 + shifted_state54_195_5 + shifted_state54_195_7);
      reservoir_sum_parallel[55] = (shifted_state55_17_0 + shifted_state55_17_1 + shifted_state55_17_3 + shifted_state55_19_2 + shifted_state55_19_4 + shifted_state55_22_0 + shifted_state55_22_4 + shifted_state55_45_1 + shifted_state55_45_2 + shifted_state55_45_4 + shifted_state55_54_1 + shifted_state55_54_3 + shifted_state55_54_5 + shifted_state55_56_1 + shifted_state55_56_4 + shifted_state55_59_1 + shifted_state55_108_0 + shifted_state55_108_1 + shifted_state55_108_2 + shifted_state55_125_2 + shifted_state55_125_3 + shifted_state55_125_5 + shifted_state55_125_7 + shifted_state55_129_0 + shifted_state55_129_2 + shifted_state55_129_3 + shifted_state55_129_5 + shifted_state55_129_6 + shifted_state55_129_7 + shifted_state55_138_0 + shifted_state55_138_1 + shifted_state55_138_2 + shifted_state55_138_3 + shifted_state55_138_4 + shifted_state55_138_5 + shifted_state55_138_6 + shifted_state55_138_7 + shifted_state55_157_2 + shifted_state55_157_4 + shifted_state55_161_1 + shifted_state55_161_3 + shifted_state55_161_6 + shifted_state55_161_7 + shifted_state55_162_0 + shifted_state55_162_2 + shifted_state55_168_0 + shifted_state55_168_1 + shifted_state55_168_4 + shifted_state55_168_5 + shifted_state55_168_6 + shifted_state55_168_7 + shifted_state55_169_2 + shifted_state55_169_4 + shifted_state55_169_5 + shifted_state55_174_0 + shifted_state55_174_5 + shifted_state55_177_2 + shifted_state55_177_3 + shifted_state55_177_4 + shifted_state55_183_5 + shifted_state55_191_1 + shifted_state55_191_2 + shifted_state55_191_3 + shifted_state55_191_4 + shifted_state55_191_6 + shifted_state55_191_7);
      reservoir_sum_parallel[56] = (shifted_state56_4_2 + shifted_state56_10_0 + shifted_state56_10_2 + shifted_state56_10_4 + shifted_state56_10_5 + shifted_state56_10_6 + shifted_state56_10_7 + shifted_state56_12_0 + shifted_state56_12_5 + shifted_state56_33_0 + shifted_state56_33_1 + shifted_state56_33_3 + shifted_state56_37_0 + shifted_state56_37_2 + shifted_state56_37_3 + shifted_state56_37_4 + shifted_state56_37_6 + shifted_state56_37_7 + shifted_state56_54_1 + shifted_state56_54_2 + shifted_state56_54_3 + shifted_state56_54_5 + shifted_state56_54_6 + shifted_state56_54_7 + shifted_state56_66_1 + shifted_state56_66_2 + shifted_state56_66_5 + shifted_state56_66_6 + shifted_state56_66_7 + shifted_state56_81_0 + shifted_state56_81_1 + shifted_state56_81_3 + shifted_state56_81_4 + shifted_state56_81_5 + shifted_state56_81_6 + shifted_state56_81_7 + shifted_state56_90_0 + shifted_state56_90_2 + shifted_state56_90_3 + shifted_state56_90_4 + shifted_state56_90_6 + shifted_state56_90_7 + shifted_state56_97_0 + shifted_state56_97_1 + shifted_state56_97_2 + shifted_state56_97_6 + shifted_state56_97_7 + shifted_state56_103_0 + shifted_state56_103_1 + shifted_state56_105_0 + shifted_state56_105_1 + shifted_state56_105_3 + shifted_state56_105_4 + shifted_state56_105_5 + shifted_state56_105_7 + shifted_state56_106_0 + shifted_state56_106_2 + shifted_state56_106_3 + shifted_state56_106_4 + shifted_state56_106_5 + shifted_state56_106_6 + shifted_state56_106_7 + shifted_state56_113_4 + shifted_state56_113_5 + shifted_state56_120_2 + shifted_state56_120_3 + shifted_state56_120_5 + shifted_state56_120_6 + shifted_state56_120_7 + shifted_state56_129_2 + shifted_state56_129_5 + shifted_state56_129_6 + shifted_state56_129_7 + shifted_state56_130_4 + shifted_state56_136_0 + shifted_state56_136_1 + shifted_state56_136_3 + shifted_state56_136_5 + shifted_state56_157_0 + shifted_state56_157_1 + shifted_state56_157_5 + shifted_state56_157_6 + shifted_state56_157_7 + shifted_state56_179_3 + shifted_state56_189_1 + shifted_state56_189_3 + shifted_state56_189_4);
      reservoir_sum_parallel[57] = (shifted_state57_34_1 + shifted_state57_34_2 + shifted_state57_34_3 + shifted_state57_34_4 + shifted_state57_34_5 + shifted_state57_34_6 + shifted_state57_34_7 + shifted_state57_51_4 + shifted_state57_55_2 + shifted_state57_55_5 + shifted_state57_58_0 + shifted_state57_58_1 + shifted_state57_58_5 + shifted_state57_58_6 + shifted_state57_58_7 + shifted_state57_78_0 + shifted_state57_78_3 + shifted_state57_78_4 + shifted_state57_78_5 + shifted_state57_78_6 + shifted_state57_78_7 + shifted_state57_104_2 + shifted_state57_104_3 + shifted_state57_105_1 + shifted_state57_105_2 + shifted_state57_105_5 + shifted_state57_115_1 + shifted_state57_115_3 + shifted_state57_137_1 + shifted_state57_137_3 + shifted_state57_137_5 + shifted_state57_142_0 + shifted_state57_142_3 + shifted_state57_142_4 + shifted_state57_147_0 + shifted_state57_147_1 + shifted_state57_147_3 + shifted_state57_147_4 + shifted_state57_154_0 + shifted_state57_154_2 + shifted_state57_154_3 + shifted_state57_154_4 + shifted_state57_154_5 + shifted_state57_154_6 + shifted_state57_154_7 + shifted_state57_156_0 + shifted_state57_156_1 + shifted_state57_156_2 + shifted_state57_156_3 + shifted_state57_156_5 + shifted_state57_164_1 + shifted_state57_164_2 + shifted_state57_164_3 + shifted_state57_164_5 + shifted_state57_164_6 + shifted_state57_164_7 + shifted_state57_167_2 + shifted_state57_167_3 + shifted_state57_167_5 + shifted_state57_167_6 + shifted_state57_167_7 + shifted_state57_173_0 + shifted_state57_173_1 + shifted_state57_173_2 + shifted_state57_173_4 + shifted_state57_177_1 + shifted_state57_177_5 + shifted_state57_177_6 + shifted_state57_177_7 + shifted_state57_179_1 + shifted_state57_179_6 + shifted_state57_179_7 + shifted_state57_181_2);
      reservoir_sum_parallel[58] = (shifted_state58_4_1 + shifted_state58_4_3 + shifted_state58_4_5 + shifted_state58_19_2 + shifted_state58_19_3 + shifted_state58_19_4 + shifted_state58_29_3 + shifted_state58_29_5 + shifted_state58_29_6 + shifted_state58_29_7 + shifted_state58_37_0 + shifted_state58_37_1 + shifted_state58_37_3 + shifted_state58_38_2 + shifted_state58_38_3 + shifted_state58_38_4 + shifted_state58_54_0 + shifted_state58_54_1 + shifted_state58_54_2 + shifted_state58_57_1 + shifted_state58_57_2 + shifted_state58_57_4 + shifted_state58_57_6 + shifted_state58_57_7 + shifted_state58_60_1 + shifted_state58_60_2 + shifted_state58_60_3 + shifted_state58_60_6 + shifted_state58_60_7 + shifted_state58_85_0 + shifted_state58_85_1 + shifted_state58_85_2 + shifted_state58_85_5 + shifted_state58_93_0 + shifted_state58_93_1 + shifted_state58_98_0 + shifted_state58_98_1 + shifted_state58_98_2 + shifted_state58_98_4 + shifted_state58_98_6 + shifted_state58_98_7 + shifted_state58_105_2 + shifted_state58_110_0 + shifted_state58_110_1 + shifted_state58_110_5 + shifted_state58_110_6 + shifted_state58_110_7 + shifted_state58_137_1 + shifted_state58_137_2 + shifted_state58_137_5 + shifted_state58_137_6 + shifted_state58_137_7 + shifted_state58_160_0 + shifted_state58_160_3 + shifted_state58_160_4 + shifted_state58_164_2 + shifted_state58_164_3 + shifted_state58_174_0 + shifted_state58_174_1 + shifted_state58_174_3 + shifted_state58_174_4 + shifted_state58_174_5 + shifted_state58_174_6 + shifted_state58_174_7);
      reservoir_sum_parallel[59] = (shifted_state59_15_0 + shifted_state59_15_1 + shifted_state59_15_2 + shifted_state59_15_3 + shifted_state59_24_0 + shifted_state59_35_0 + shifted_state59_35_1 + shifted_state59_35_2 + shifted_state59_35_5 + shifted_state59_44_0 + shifted_state59_44_3 + shifted_state59_44_5 + shifted_state59_44_6 + shifted_state59_44_7 + shifted_state59_46_1 + shifted_state59_46_4 + shifted_state59_47_0 + shifted_state59_90_3 + shifted_state59_90_4 + shifted_state59_90_6 + shifted_state59_90_7 + shifted_state59_98_2 + shifted_state59_98_3 + shifted_state59_105_1 + shifted_state59_105_2 + shifted_state59_105_3 + shifted_state59_105_5 + shifted_state59_105_6 + shifted_state59_105_7 + shifted_state59_115_0 + shifted_state59_115_1 + shifted_state59_115_2 + shifted_state59_115_4 + shifted_state59_115_5 + shifted_state59_115_6 + shifted_state59_115_7 + shifted_state59_116_2 + shifted_state59_116_3 + shifted_state59_116_5 + shifted_state59_121_3 + shifted_state59_121_4 + shifted_state59_121_5 + shifted_state59_121_6 + shifted_state59_121_7 + shifted_state59_136_0 + shifted_state59_136_1 + shifted_state59_136_2 + shifted_state59_136_3 + shifted_state59_136_5 + shifted_state59_138_0 + shifted_state59_138_5 + shifted_state59_138_6 + shifted_state59_138_7 + shifted_state59_157_2 + shifted_state59_157_4 + shifted_state59_157_5 + shifted_state59_180_0 + shifted_state59_180_1 + shifted_state59_180_5 + shifted_state59_180_6 + shifted_state59_180_7 + shifted_state59_194_1 + shifted_state59_194_4 + shifted_state59_194_6 + shifted_state59_194_7 + shifted_state59_198_3 + shifted_state59_198_4 + shifted_state59_198_5 + shifted_state59_198_6 + shifted_state59_198_7);
      reservoir_sum_parallel[60] = (shifted_state60_3_2 + shifted_state60_10_0 + shifted_state60_10_1 + shifted_state60_10_4 + shifted_state60_10_5 + shifted_state60_10_6 + shifted_state60_10_7 + shifted_state60_20_0 + shifted_state60_20_1 + shifted_state60_20_2 + shifted_state60_20_4 + shifted_state60_20_5 + shifted_state60_20_6 + shifted_state60_20_7 + shifted_state60_24_0 + shifted_state60_24_1 + shifted_state60_24_2 + shifted_state60_24_3 + shifted_state60_24_4 + shifted_state60_28_0 + shifted_state60_28_1 + shifted_state60_28_2 + shifted_state60_28_4 + shifted_state60_46_2 + shifted_state60_46_5 + shifted_state60_46_6 + shifted_state60_46_7 + shifted_state60_63_0 + shifted_state60_63_1 + shifted_state60_63_2 + shifted_state60_63_3 + shifted_state60_63_5 + shifted_state60_63_6 + shifted_state60_63_7 + shifted_state60_72_5 + shifted_state60_84_0 + shifted_state60_91_0 + shifted_state60_91_5 + shifted_state60_91_6 + shifted_state60_91_7 + shifted_state60_109_0 + shifted_state60_109_2 + shifted_state60_109_3 + shifted_state60_109_4 + shifted_state60_109_5 + shifted_state60_109_6 + shifted_state60_109_7 + shifted_state60_116_1 + shifted_state60_116_3 + shifted_state60_123_0 + shifted_state60_123_1 + shifted_state60_123_3 + shifted_state60_123_5 + shifted_state60_125_0 + shifted_state60_125_3 + shifted_state60_137_0 + shifted_state60_137_3 + shifted_state60_137_4 + shifted_state60_137_5 + shifted_state60_137_6 + shifted_state60_137_7 + shifted_state60_139_0 + shifted_state60_139_1 + shifted_state60_139_2 + shifted_state60_139_4 + shifted_state60_169_0 + shifted_state60_169_3 + shifted_state60_169_4 + shifted_state60_169_6 + shifted_state60_169_7 + shifted_state60_170_0 + shifted_state60_170_1 + shifted_state60_170_3 + shifted_state60_170_6 + shifted_state60_177_0 + shifted_state60_177_1 + shifted_state60_177_2 + shifted_state60_177_3 + shifted_state60_177_4 + shifted_state60_177_6 + shifted_state60_177_7 + shifted_state60_195_0 + shifted_state60_195_3);
      reservoir_sum_parallel[61] = (shifted_state61_1_0 + shifted_state61_1_2 + shifted_state61_1_4 + shifted_state61_5_0 + shifted_state61_5_3 + shifted_state61_11_0 + shifted_state61_11_4 + shifted_state61_14_2 + shifted_state61_31_3 + shifted_state61_31_4 + shifted_state61_34_0 + shifted_state61_34_3 + shifted_state61_34_4 + shifted_state61_34_6 + shifted_state61_34_7 + shifted_state61_35_0 + shifted_state61_35_1 + shifted_state61_35_2 + shifted_state61_35_4 + shifted_state61_50_0 + shifted_state61_50_1 + shifted_state61_50_6 + shifted_state61_59_0 + shifted_state61_59_4 + shifted_state61_59_5 + shifted_state61_59_6 + shifted_state61_59_7 + shifted_state61_84_3 + shifted_state61_84_5 + shifted_state61_86_0 + shifted_state61_86_2 + shifted_state61_86_4 + shifted_state61_86_6 + shifted_state61_86_7 + shifted_state61_89_0 + shifted_state61_89_2 + shifted_state61_95_0 + shifted_state61_95_1 + shifted_state61_95_4 + shifted_state61_99_3 + shifted_state61_99_4 + shifted_state61_117_2 + shifted_state61_117_4 + shifted_state61_117_5 + shifted_state61_118_1 + shifted_state61_118_4 + shifted_state61_118_5 + shifted_state61_118_6 + shifted_state61_118_7 + shifted_state61_119_0 + shifted_state61_119_5 + shifted_state61_119_6 + shifted_state61_119_7 + shifted_state61_122_3 + shifted_state61_122_4 + shifted_state61_122_5 + shifted_state61_122_6 + shifted_state61_122_7 + shifted_state61_123_0 + shifted_state61_123_1 + shifted_state61_123_2 + shifted_state61_123_4 + shifted_state61_134_1 + shifted_state61_134_3 + shifted_state61_136_5 + shifted_state61_136_6 + shifted_state61_136_7 + shifted_state61_142_0 + shifted_state61_142_1 + shifted_state61_142_5 + shifted_state61_142_6 + shifted_state61_142_7 + shifted_state61_148_0 + shifted_state61_148_1 + shifted_state61_148_5 + shifted_state61_152_0 + shifted_state61_152_1 + shifted_state61_152_2 + shifted_state61_152_3 + shifted_state61_163_0 + shifted_state61_163_2 + shifted_state61_163_3 + shifted_state61_163_5 + shifted_state61_163_6 + shifted_state61_163_7 + shifted_state61_164_2 + shifted_state61_175_3 + shifted_state61_179_4 + shifted_state61_179_5);
      reservoir_sum_parallel[62] = (shifted_state62_9_0 + shifted_state62_9_2 + shifted_state62_14_0 + shifted_state62_14_3 + shifted_state62_14_4 + shifted_state62_14_5 + shifted_state62_14_6 + shifted_state62_14_7 + shifted_state62_19_0 + shifted_state62_19_2 + shifted_state62_19_3 + shifted_state62_19_4 + shifted_state62_29_0 + shifted_state62_29_1 + shifted_state62_29_4 + shifted_state62_35_1 + shifted_state62_35_2 + shifted_state62_47_2 + shifted_state62_47_3 + shifted_state62_47_5 + shifted_state62_47_6 + shifted_state62_47_7 + shifted_state62_67_0 + shifted_state62_67_1 + shifted_state62_67_2 + shifted_state62_67_5 + shifted_state62_107_0 + shifted_state62_107_1 + shifted_state62_121_0 + shifted_state62_121_1 + shifted_state62_121_2 + shifted_state62_121_4 + shifted_state62_130_2 + shifted_state62_130_4 + shifted_state62_130_6 + shifted_state62_130_7 + shifted_state62_134_0 + shifted_state62_134_1 + shifted_state62_134_5 + shifted_state62_134_6 + shifted_state62_134_7 + shifted_state62_137_1 + shifted_state62_137_3 + shifted_state62_137_6 + shifted_state62_137_7 + shifted_state62_138_0 + shifted_state62_138_5 + shifted_state62_143_0 + shifted_state62_143_2 + shifted_state62_143_4 + shifted_state62_162_0 + shifted_state62_162_2 + shifted_state62_178_0 + shifted_state62_178_2 + shifted_state62_178_3 + shifted_state62_178_4 + shifted_state62_178_5 + shifted_state62_178_6 + shifted_state62_178_7 + shifted_state62_181_2 + shifted_state62_181_4 + shifted_state62_181_6 + shifted_state62_181_7 + shifted_state62_189_3 + shifted_state62_189_5 + shifted_state62_189_6 + shifted_state62_189_7);
      reservoir_sum_parallel[63] = (shifted_state63_4_2 + shifted_state63_4_3 + shifted_state63_11_0 + shifted_state63_11_1 + shifted_state63_11_3 + shifted_state63_11_4 + shifted_state63_11_5 + shifted_state63_11_6 + shifted_state63_11_7 + shifted_state63_37_0 + shifted_state63_37_4 + shifted_state63_37_5 + shifted_state63_37_6 + shifted_state63_37_7 + shifted_state63_43_0 + shifted_state63_43_1 + shifted_state63_43_3 + shifted_state63_43_4 + shifted_state63_43_5 + shifted_state63_43_6 + shifted_state63_43_7 + shifted_state63_73_5 + shifted_state63_73_6 + shifted_state63_73_7 + shifted_state63_87_4 + shifted_state63_89_1 + shifted_state63_89_3 + shifted_state63_89_4 + shifted_state63_91_0 + shifted_state63_91_3 + shifted_state63_91_5 + shifted_state63_91_6 + shifted_state63_91_7 + shifted_state63_92_0 + shifted_state63_92_2 + shifted_state63_92_3 + shifted_state63_92_5 + shifted_state63_92_6 + shifted_state63_92_7 + shifted_state63_100_0 + shifted_state63_100_1 + shifted_state63_100_6 + shifted_state63_100_7 + shifted_state63_104_1 + shifted_state63_104_2 + shifted_state63_104_3 + shifted_state63_104_5 + shifted_state63_104_6 + shifted_state63_104_7 + shifted_state63_127_0 + shifted_state63_127_1 + shifted_state63_127_2 + shifted_state63_127_3 + shifted_state63_128_0 + shifted_state63_128_1 + shifted_state63_128_2 + shifted_state63_129_0 + shifted_state63_129_6 + shifted_state63_129_7 + shifted_state63_131_1 + shifted_state63_131_2 + shifted_state63_131_3 + shifted_state63_131_6 + shifted_state63_131_7 + shifted_state63_138_0 + shifted_state63_138_2 + shifted_state63_138_3 + shifted_state63_138_5 + shifted_state63_138_6 + shifted_state63_138_7 + shifted_state63_155_2 + shifted_state63_155_3 + shifted_state63_155_6 + shifted_state63_165_1 + shifted_state63_165_3 + shifted_state63_165_5 + shifted_state63_184_0 + shifted_state63_184_4 + shifted_state63_184_6 + shifted_state63_184_7 + shifted_state63_195_0 + shifted_state63_195_1 + shifted_state63_195_3 + shifted_state63_195_5 + shifted_state63_195_6 + shifted_state63_195_7);
      reservoir_sum_parallel[64] = (shifted_state64_23_1 + shifted_state64_23_2 + shifted_state64_23_3 + shifted_state64_26_1 + shifted_state64_26_2 + shifted_state64_26_3 + shifted_state64_26_4 + shifted_state64_26_5 + shifted_state64_26_6 + shifted_state64_26_7 + shifted_state64_30_0 + shifted_state64_30_1 + shifted_state64_38_1 + shifted_state64_38_2 + shifted_state64_38_3 + shifted_state64_64_0 + shifted_state64_64_1 + shifted_state64_65_1 + shifted_state64_83_0 + shifted_state64_83_1 + shifted_state64_83_2 + shifted_state64_83_3 + shifted_state64_92_2 + shifted_state64_92_5 + shifted_state64_93_0 + shifted_state64_93_1 + shifted_state64_93_2 + shifted_state64_93_5 + shifted_state64_93_6 + shifted_state64_93_7 + shifted_state64_98_0 + shifted_state64_98_1 + shifted_state64_98_4 + shifted_state64_98_6 + shifted_state64_98_7 + shifted_state64_103_0 + shifted_state64_103_2 + shifted_state64_103_4 + shifted_state64_103_5 + shifted_state64_103_6 + shifted_state64_103_7 + shifted_state64_122_0 + shifted_state64_122_2 + shifted_state64_122_4 + shifted_state64_123_0 + shifted_state64_123_1 + shifted_state64_123_2 + shifted_state64_123_3 + shifted_state64_123_4 + shifted_state64_123_5 + shifted_state64_123_6 + shifted_state64_123_7 + shifted_state64_128_0 + shifted_state64_128_1 + shifted_state64_128_3 + shifted_state64_131_1 + shifted_state64_131_3 + shifted_state64_131_5 + shifted_state64_131_6 + shifted_state64_131_7 + shifted_state64_134_0 + shifted_state64_134_1 + shifted_state64_134_3 + shifted_state64_134_4 + shifted_state64_134_6 + shifted_state64_134_7 + shifted_state64_174_1 + shifted_state64_174_3 + shifted_state64_174_5 + shifted_state64_174_6 + shifted_state64_174_7 + shifted_state64_177_0 + shifted_state64_177_1 + shifted_state64_177_3 + shifted_state64_177_6 + shifted_state64_177_7 + shifted_state64_181_0 + shifted_state64_181_3 + shifted_state64_181_4 + shifted_state64_181_5 + shifted_state64_181_6 + shifted_state64_181_7 + shifted_state64_184_0 + shifted_state64_184_3 + shifted_state64_184_5 + shifted_state64_188_0 + shifted_state64_188_1 + shifted_state64_188_2);
      reservoir_sum_parallel[65] = (shifted_state65_3_0 + shifted_state65_3_5 + shifted_state65_3_6 + shifted_state65_3_7 + shifted_state65_10_0 + shifted_state65_10_2 + shifted_state65_10_3 + shifted_state65_10_6 + shifted_state65_10_7 + shifted_state65_11_0 + shifted_state65_11_3 + shifted_state65_11_4 + shifted_state65_11_5 + shifted_state65_11_6 + shifted_state65_11_7 + shifted_state65_13_1 + shifted_state65_13_3 + shifted_state65_13_4 + shifted_state65_19_0 + shifted_state65_19_3 + shifted_state65_19_4 + shifted_state65_19_5 + shifted_state65_19_6 + shifted_state65_19_7 + shifted_state65_21_0 + shifted_state65_21_5 + shifted_state65_64_1 + shifted_state65_64_2 + shifted_state65_64_3 + shifted_state65_96_1 + shifted_state65_96_2 + shifted_state65_96_3 + shifted_state65_96_5 + shifted_state65_99_0 + shifted_state65_99_1 + shifted_state65_99_5 + shifted_state65_110_0 + shifted_state65_110_5 + shifted_state65_111_0 + shifted_state65_111_3 + shifted_state65_111_4 + shifted_state65_111_5 + shifted_state65_111_6 + shifted_state65_111_7 + shifted_state65_119_1 + shifted_state65_119_2 + shifted_state65_136_4 + shifted_state65_146_3 + shifted_state65_146_4 + shifted_state65_152_0 + shifted_state65_152_1 + shifted_state65_152_2 + shifted_state65_152_3 + shifted_state65_152_4 + shifted_state65_152_5 + shifted_state65_152_6 + shifted_state65_152_7 + shifted_state65_156_0 + shifted_state65_165_0 + shifted_state65_165_1 + shifted_state65_165_2 + shifted_state65_174_1 + shifted_state65_174_3 + shifted_state65_182_0 + shifted_state65_182_2 + shifted_state65_182_5 + shifted_state65_188_0 + shifted_state65_188_3 + shifted_state65_188_4);
      reservoir_sum_parallel[66] = (shifted_state66_7_0 + shifted_state66_7_1 + shifted_state66_7_3 + shifted_state66_15_0 + shifted_state66_15_1 + shifted_state66_15_2 + shifted_state66_15_4 + shifted_state66_15_6 + shifted_state66_15_7 + shifted_state66_22_0 + shifted_state66_22_1 + shifted_state66_22_3 + shifted_state66_28_1 + shifted_state66_28_2 + shifted_state66_28_5 + shifted_state66_28_6 + shifted_state66_28_7 + shifted_state66_61_1 + shifted_state66_61_2 + shifted_state66_61_5 + shifted_state66_96_1 + shifted_state66_96_5 + shifted_state66_99_4 + shifted_state66_99_5 + shifted_state66_99_6 + shifted_state66_99_7 + shifted_state66_103_5 + shifted_state66_103_6 + shifted_state66_103_7 + shifted_state66_107_0 + shifted_state66_107_1 + shifted_state66_107_2 + shifted_state66_107_3 + shifted_state66_107_5 + shifted_state66_107_6 + shifted_state66_107_7 + shifted_state66_112_2 + shifted_state66_112_6 + shifted_state66_112_7 + shifted_state66_115_4 + shifted_state66_117_0 + shifted_state66_117_1 + shifted_state66_117_2 + shifted_state66_117_3 + shifted_state66_119_0 + shifted_state66_119_4 + shifted_state66_127_3 + shifted_state66_127_6 + shifted_state66_127_7 + shifted_state66_163_1 + shifted_state66_163_2 + shifted_state66_163_3 + shifted_state66_163_4 + shifted_state66_168_0 + shifted_state66_168_2 + shifted_state66_168_3 + shifted_state66_168_5 + shifted_state66_168_6 + shifted_state66_168_7 + shifted_state66_189_0 + shifted_state66_189_3 + shifted_state66_192_2);
      reservoir_sum_parallel[67] = (shifted_state67_0_1 + shifted_state67_0_3 + shifted_state67_0_4 + shifted_state67_0_6 + shifted_state67_0_7 + shifted_state67_5_2 + shifted_state67_5_3 + shifted_state67_5_4 + shifted_state67_5_5 + shifted_state67_28_0 + shifted_state67_28_5 + shifted_state67_28_6 + shifted_state67_28_7 + shifted_state67_31_0 + shifted_state67_31_2 + shifted_state67_33_0 + shifted_state67_55_0 + shifted_state67_55_1 + shifted_state67_55_3 + shifted_state67_55_5 + shifted_state67_55_6 + shifted_state67_55_7 + shifted_state67_61_0 + shifted_state67_61_1 + shifted_state67_61_3 + shifted_state67_61_4 + shifted_state67_61_5 + shifted_state67_61_6 + shifted_state67_61_7 + shifted_state67_64_0 + shifted_state67_64_1 + shifted_state67_64_2 + shifted_state67_64_3 + shifted_state67_64_4 + shifted_state67_64_5 + shifted_state67_64_6 + shifted_state67_64_7 + shifted_state67_86_3 + shifted_state67_86_5 + shifted_state67_86_6 + shifted_state67_86_7 + shifted_state67_90_0 + shifted_state67_90_1 + shifted_state67_90_2 + shifted_state67_90_5 + shifted_state67_90_6 + shifted_state67_90_7 + shifted_state67_120_3 + shifted_state67_120_6 + shifted_state67_133_0 + shifted_state67_133_1 + shifted_state67_133_3 + shifted_state67_133_4 + shifted_state67_144_1 + shifted_state67_144_2 + shifted_state67_144_4 + shifted_state67_156_0 + shifted_state67_156_1 + shifted_state67_156_2 + shifted_state67_165_0 + shifted_state67_165_1 + shifted_state67_165_3 + shifted_state67_165_4 + shifted_state67_165_5 + shifted_state67_165_6 + shifted_state67_165_7 + shifted_state67_170_0 + shifted_state67_170_1 + shifted_state67_190_0 + shifted_state67_190_1 + shifted_state67_190_2 + shifted_state67_190_4 + shifted_state67_190_6 + shifted_state67_190_7);
      reservoir_sum_parallel[68] = (shifted_state68_8_1 + shifted_state68_8_3 + shifted_state68_23_1 + shifted_state68_23_2 + shifted_state68_23_3 + shifted_state68_23_5 + shifted_state68_23_6 + shifted_state68_23_7 + shifted_state68_29_4 + shifted_state68_36_0 + shifted_state68_36_3 + shifted_state68_53_5 + shifted_state68_53_6 + shifted_state68_53_7 + shifted_state68_61_2 + shifted_state68_61_3 + shifted_state68_61_4 + shifted_state68_61_5 + shifted_state68_61_6 + shifted_state68_61_7 + shifted_state68_91_2 + shifted_state68_95_0 + shifted_state68_95_1 + shifted_state68_95_3 + shifted_state68_95_4 + shifted_state68_95_5 + shifted_state68_95_6 + shifted_state68_95_7 + shifted_state68_106_2 + shifted_state68_106_4 + shifted_state68_106_6 + shifted_state68_106_7 + shifted_state68_107_1 + shifted_state68_107_2 + shifted_state68_107_3 + shifted_state68_107_4 + shifted_state68_107_5 + shifted_state68_107_6 + shifted_state68_107_7 + shifted_state68_121_1 + shifted_state68_121_5 + shifted_state68_125_3 + shifted_state68_133_0 + shifted_state68_133_1 + shifted_state68_133_3 + shifted_state68_133_4 + shifted_state68_133_6 + shifted_state68_133_7 + shifted_state68_148_0 + shifted_state68_148_2 + shifted_state68_148_3 + shifted_state68_148_5 + shifted_state68_148_6 + shifted_state68_148_7 + shifted_state68_152_1 + shifted_state68_152_2 + shifted_state68_152_4 + shifted_state68_152_5 + shifted_state68_152_6 + shifted_state68_152_7 + shifted_state68_159_2 + shifted_state68_159_3 + shifted_state68_159_4 + shifted_state68_159_6 + shifted_state68_159_7 + shifted_state68_175_0 + shifted_state68_175_2 + shifted_state68_175_3 + shifted_state68_175_6 + shifted_state68_175_7 + shifted_state68_182_3 + shifted_state68_182_5);
      reservoir_sum_parallel[69] = (shifted_state69_2_1 + shifted_state69_2_2 + shifted_state69_2_4 + shifted_state69_2_5 + shifted_state69_2_6 + shifted_state69_2_7 + shifted_state69_26_1 + shifted_state69_26_3 + shifted_state69_26_5 + shifted_state69_26_6 + shifted_state69_26_7 + shifted_state69_34_0 + shifted_state69_34_3 + shifted_state69_34_4 + shifted_state69_34_5 + shifted_state69_34_6 + shifted_state69_34_7 + shifted_state69_36_0 + shifted_state69_36_3 + shifted_state69_46_0 + shifted_state69_46_2 + shifted_state69_46_3 + shifted_state69_46_4 + shifted_state69_46_5 + shifted_state69_46_6 + shifted_state69_46_7 + shifted_state69_49_0 + shifted_state69_49_3 + shifted_state69_49_5 + shifted_state69_52_3 + shifted_state69_64_0 + shifted_state69_64_1 + shifted_state69_64_2 + shifted_state69_64_4 + shifted_state69_64_6 + shifted_state69_64_7 + shifted_state69_74_0 + shifted_state69_74_1 + shifted_state69_93_2 + shifted_state69_93_3 + shifted_state69_93_5 + shifted_state69_93_6 + shifted_state69_93_7 + shifted_state69_100_0 + shifted_state69_100_3 + shifted_state69_109_0 + shifted_state69_109_5 + shifted_state69_109_6 + shifted_state69_109_7 + shifted_state69_111_0 + shifted_state69_111_1 + shifted_state69_111_3 + shifted_state69_111_4 + shifted_state69_111_5 + shifted_state69_111_6 + shifted_state69_111_7 + shifted_state69_132_2 + shifted_state69_132_3 + shifted_state69_132_4 + shifted_state69_132_5 + shifted_state69_148_1 + shifted_state69_148_3 + shifted_state69_148_5 + shifted_state69_148_6 + shifted_state69_148_7 + shifted_state69_175_0 + shifted_state69_175_1 + shifted_state69_175_2 + shifted_state69_175_3 + shifted_state69_175_4 + shifted_state69_175_6 + shifted_state69_175_7 + shifted_state69_183_0 + shifted_state69_183_2);
      reservoir_sum_parallel[70] = (shifted_state70_1_4 + shifted_state70_28_1 + shifted_state70_28_2 + shifted_state70_28_3 + shifted_state70_43_2 + shifted_state70_43_3 + shifted_state70_43_5 + shifted_state70_66_1 + shifted_state70_66_6 + shifted_state70_66_7 + shifted_state70_105_0 + shifted_state70_105_1 + shifted_state70_105_5 + shifted_state70_118_0 + shifted_state70_118_3 + shifted_state70_118_4 + shifted_state70_126_0 + shifted_state70_126_2 + shifted_state70_126_3 + shifted_state70_126_4 + shifted_state70_126_5 + shifted_state70_126_6 + shifted_state70_126_7 + shifted_state70_128_0 + shifted_state70_128_2 + shifted_state70_128_5 + shifted_state70_128_6 + shifted_state70_128_7 + shifted_state70_155_0 + shifted_state70_155_1 + shifted_state70_158_1 + shifted_state70_162_0 + shifted_state70_162_2 + shifted_state70_162_5 + shifted_state70_162_6 + shifted_state70_162_7 + shifted_state70_165_1 + shifted_state70_165_2 + shifted_state70_182_0 + shifted_state70_182_1 + shifted_state70_182_2 + shifted_state70_182_4 + shifted_state70_182_5 + shifted_state70_182_6 + shifted_state70_182_7 + shifted_state70_188_0 + shifted_state70_188_1 + shifted_state70_188_2 + shifted_state70_188_3 + shifted_state70_188_4 + shifted_state70_188_5 + shifted_state70_188_6 + shifted_state70_188_7);
      reservoir_sum_parallel[71] = (shifted_state71_13_0 + shifted_state71_13_2 + shifted_state71_39_1 + shifted_state71_39_4 + shifted_state71_39_5 + shifted_state71_39_6 + shifted_state71_39_7 + shifted_state71_47_2 + shifted_state71_47_3 + shifted_state71_47_4 + shifted_state71_47_5 + shifted_state71_47_6 + shifted_state71_47_7 + shifted_state71_61_0 + shifted_state71_61_2 + shifted_state71_61_6 + shifted_state71_61_7 + shifted_state71_90_0 + shifted_state71_90_2 + shifted_state71_90_3 + shifted_state71_90_5 + shifted_state71_90_6 + shifted_state71_90_7 + shifted_state71_96_0 + shifted_state71_96_3 + shifted_state71_96_4 + shifted_state71_96_6 + shifted_state71_96_7 + shifted_state71_103_0 + shifted_state71_103_2 + shifted_state71_103_3 + shifted_state71_104_1 + shifted_state71_104_5 + shifted_state71_151_0 + shifted_state71_151_1 + shifted_state71_151_3 + shifted_state71_151_4 + shifted_state71_151_5 + shifted_state71_151_7 + shifted_state71_153_2 + shifted_state71_155_0 + shifted_state71_155_1 + shifted_state71_155_2 + shifted_state71_155_3 + shifted_state71_155_6 + shifted_state71_155_7 + shifted_state71_169_0 + shifted_state71_169_1 + shifted_state71_169_4 + shifted_state71_169_5 + shifted_state71_169_6 + shifted_state71_169_7 + shifted_state71_173_0 + shifted_state71_173_2 + shifted_state71_173_3 + shifted_state71_173_4);
      reservoir_sum_parallel[72] = (shifted_state72_2_0 + shifted_state72_2_4 + shifted_state72_20_0 + shifted_state72_20_2 + shifted_state72_20_6 + shifted_state72_22_1 + shifted_state72_22_3 + shifted_state72_25_0 + shifted_state72_25_1 + shifted_state72_25_2 + shifted_state72_25_3 + shifted_state72_25_5 + shifted_state72_26_1 + shifted_state72_26_3 + shifted_state72_26_4 + shifted_state72_35_2 + shifted_state72_35_4 + shifted_state72_35_6 + shifted_state72_35_7 + shifted_state72_38_4 + shifted_state72_38_5 + shifted_state72_38_6 + shifted_state72_38_7 + shifted_state72_66_0 + shifted_state72_66_1 + shifted_state72_66_3 + shifted_state72_68_0 + shifted_state72_68_3 + shifted_state72_68_4 + shifted_state72_69_0 + shifted_state72_69_1 + shifted_state72_69_3 + shifted_state72_70_3 + shifted_state72_70_5 + shifted_state72_70_6 + shifted_state72_70_7 + shifted_state72_79_0 + shifted_state72_79_3 + shifted_state72_79_4 + shifted_state72_79_6 + shifted_state72_79_7 + shifted_state72_86_6 + shifted_state72_102_0 + shifted_state72_102_1 + shifted_state72_102_2 + shifted_state72_102_3 + shifted_state72_109_1 + shifted_state72_109_3 + shifted_state72_109_4 + shifted_state72_111_0 + shifted_state72_111_1 + shifted_state72_111_2 + shifted_state72_125_0 + shifted_state72_125_1 + shifted_state72_125_3 + shifted_state72_125_4 + shifted_state72_125_5 + shifted_state72_125_6 + shifted_state72_125_7 + shifted_state72_137_0 + shifted_state72_137_1 + shifted_state72_137_3 + shifted_state72_137_4 + shifted_state72_137_5 + shifted_state72_137_6 + shifted_state72_137_7 + shifted_state72_143_0 + shifted_state72_143_1 + shifted_state72_143_3 + shifted_state72_143_4 + shifted_state72_143_5 + shifted_state72_143_6 + shifted_state72_143_7 + shifted_state72_144_0 + shifted_state72_144_2 + shifted_state72_144_3 + shifted_state72_152_0 + shifted_state72_152_4 + shifted_state72_152_5 + shifted_state72_152_7 + shifted_state72_177_0 + shifted_state72_177_1 + shifted_state72_177_2 + shifted_state72_177_5 + shifted_state72_177_6 + shifted_state72_177_7 + shifted_state72_178_0 + shifted_state72_178_1 + shifted_state72_186_1 + shifted_state72_186_2 + shifted_state72_186_3);
      reservoir_sum_parallel[73] = (shifted_state73_5_1 + shifted_state73_5_3 + shifted_state73_42_1 + shifted_state73_42_3 + shifted_state73_42_4 + shifted_state73_42_5 + shifted_state73_43_1 + shifted_state73_43_3 + shifted_state73_43_4 + shifted_state73_43_5 + shifted_state73_43_6 + shifted_state73_43_7 + shifted_state73_52_0 + shifted_state73_52_3 + shifted_state73_70_2 + shifted_state73_70_4 + shifted_state73_70_5 + shifted_state73_70_6 + shifted_state73_70_7 + shifted_state73_72_0 + shifted_state73_72_2 + shifted_state73_72_3 + shifted_state73_72_4 + shifted_state73_72_6 + shifted_state73_72_7 + shifted_state73_110_0 + shifted_state73_110_2 + shifted_state73_110_5 + shifted_state73_111_0 + shifted_state73_111_1 + shifted_state73_111_3 + shifted_state73_114_0 + shifted_state73_114_1 + shifted_state73_114_2 + shifted_state73_114_3 + shifted_state73_114_6 + shifted_state73_114_7 + shifted_state73_123_0 + shifted_state73_123_2 + shifted_state73_123_4 + shifted_state73_123_5 + shifted_state73_123_6 + shifted_state73_123_7 + shifted_state73_129_0 + shifted_state73_129_2 + shifted_state73_129_3 + shifted_state73_129_4 + shifted_state73_138_1 + shifted_state73_138_4 + shifted_state73_138_5 + shifted_state73_138_6 + shifted_state73_138_7 + shifted_state73_150_2 + shifted_state73_150_5 + shifted_state73_150_6 + shifted_state73_150_7 + shifted_state73_164_0 + shifted_state73_164_1 + shifted_state73_164_2 + shifted_state73_177_0 + shifted_state73_177_3 + shifted_state73_177_5 + shifted_state73_177_6 + shifted_state73_177_7 + shifted_state73_179_0 + shifted_state73_179_4 + shifted_state73_180_0 + shifted_state73_180_1 + shifted_state73_180_2 + shifted_state73_180_4 + shifted_state73_181_0 + shifted_state73_181_2 + shifted_state73_181_5 + shifted_state73_182_0 + shifted_state73_182_2 + shifted_state73_182_4 + shifted_state73_182_5 + shifted_state73_182_7 + shifted_state73_193_1 + shifted_state73_193_3 + shifted_state73_193_4 + shifted_state73_193_5 + shifted_state73_195_0 + shifted_state73_195_1 + shifted_state73_195_4 + shifted_state73_195_5 + shifted_state73_195_6 + shifted_state73_195_7);
      reservoir_sum_parallel[74] = (shifted_state74_6_1 + shifted_state74_6_2 + shifted_state74_6_3 + shifted_state74_13_1 + shifted_state74_13_3 + shifted_state74_13_4 + shifted_state74_13_5 + shifted_state74_13_6 + shifted_state74_13_7 + shifted_state74_16_0 + shifted_state74_16_5 + shifted_state74_16_6 + shifted_state74_16_7 + shifted_state74_24_0 + shifted_state74_24_1 + shifted_state74_24_2 + shifted_state74_24_3 + shifted_state74_24_4 + shifted_state74_24_5 + shifted_state74_24_6 + shifted_state74_24_7 + shifted_state74_31_0 + shifted_state74_31_1 + shifted_state74_31_4 + shifted_state74_31_5 + shifted_state74_55_1 + shifted_state74_55_4 + shifted_state74_55_5 + shifted_state74_55_6 + shifted_state74_55_7 + shifted_state74_81_3 + shifted_state74_81_4 + shifted_state74_83_0 + shifted_state74_83_1 + shifted_state74_83_3 + shifted_state74_83_4 + shifted_state74_83_5 + shifted_state74_83_6 + shifted_state74_83_7 + shifted_state74_85_0 + shifted_state74_85_1 + shifted_state74_85_4 + shifted_state74_85_5 + shifted_state74_85_6 + shifted_state74_85_7 + shifted_state74_89_0 + shifted_state74_89_1 + shifted_state74_89_2 + shifted_state74_89_3 + shifted_state74_89_4 + shifted_state74_89_5 + shifted_state74_89_6 + shifted_state74_89_7 + shifted_state74_95_1 + shifted_state74_95_2 + shifted_state74_95_3 + shifted_state74_95_4 + shifted_state74_98_0 + shifted_state74_98_1 + shifted_state74_98_2 + shifted_state74_98_3 + shifted_state74_98_5 + shifted_state74_98_7 + shifted_state74_118_0 + shifted_state74_118_2 + shifted_state74_118_3 + shifted_state74_118_4 + shifted_state74_118_5 + shifted_state74_118_6 + shifted_state74_118_7 + shifted_state74_121_0 + shifted_state74_121_1 + shifted_state74_121_3 + shifted_state74_121_4 + shifted_state74_121_5 + shifted_state74_121_7 + shifted_state74_123_1 + shifted_state74_123_3 + shifted_state74_126_0 + shifted_state74_126_2 + shifted_state74_126_4 + shifted_state74_138_0 + shifted_state74_138_1 + shifted_state74_138_4 + shifted_state74_138_6 + shifted_state74_138_7 + shifted_state74_149_0 + shifted_state74_149_2 + shifted_state74_149_4 + shifted_state74_150_0 + shifted_state74_150_1 + shifted_state74_150_2 + shifted_state74_157_3 + shifted_state74_157_4 + shifted_state74_157_6 + shifted_state74_157_7 + shifted_state74_166_2 + shifted_state74_166_4 + shifted_state74_176_0 + shifted_state74_176_1 + shifted_state74_176_3 + shifted_state74_176_5 + shifted_state74_176_6 + shifted_state74_176_7 + shifted_state74_194_2 + shifted_state74_194_3 + shifted_state74_194_4 + shifted_state74_194_5);
      reservoir_sum_parallel[75] = (shifted_state75_14_4 + shifted_state75_14_5 + shifted_state75_14_6 + shifted_state75_14_7 + shifted_state75_38_0 + shifted_state75_38_3 + shifted_state75_38_5 + shifted_state75_42_1 + shifted_state75_42_2 + shifted_state75_42_3 + shifted_state75_42_4 + shifted_state75_42_6 + shifted_state75_42_7 + shifted_state75_53_1 + shifted_state75_53_4 + shifted_state75_53_5 + shifted_state75_53_6 + shifted_state75_53_7 + shifted_state75_56_2 + shifted_state75_56_3 + shifted_state75_65_1 + shifted_state75_86_1 + shifted_state75_86_4 + shifted_state75_88_4 + shifted_state75_88_5 + shifted_state75_88_6 + shifted_state75_88_7 + shifted_state75_93_1 + shifted_state75_93_2 + shifted_state75_93_6 + shifted_state75_93_7 + shifted_state75_99_0 + shifted_state75_99_2 + shifted_state75_99_5 + shifted_state75_100_1 + shifted_state75_100_5 + shifted_state75_105_1 + shifted_state75_105_2 + shifted_state75_105_3 + shifted_state75_105_4 + shifted_state75_105_5 + shifted_state75_105_6 + shifted_state75_105_7 + shifted_state75_108_0 + shifted_state75_108_1 + shifted_state75_108_4 + shifted_state75_108_5 + shifted_state75_108_6 + shifted_state75_108_7 + shifted_state75_126_2 + shifted_state75_126_3 + shifted_state75_126_5 + shifted_state75_126_6 + shifted_state75_126_7 + shifted_state75_131_0 + shifted_state75_131_5 + shifted_state75_134_2 + shifted_state75_134_5 + shifted_state75_146_0 + shifted_state75_146_1 + shifted_state75_146_3 + shifted_state75_146_5 + shifted_state75_146_6 + shifted_state75_146_7 + shifted_state75_151_0 + shifted_state75_151_1 + shifted_state75_151_3 + shifted_state75_151_5 + shifted_state75_151_6 + shifted_state75_151_7 + shifted_state75_164_4 + shifted_state75_167_1 + shifted_state75_167_2 + shifted_state75_169_4 + shifted_state75_169_5 + shifted_state75_182_0 + shifted_state75_182_4 + shifted_state75_182_5 + shifted_state75_182_6 + shifted_state75_182_7 + shifted_state75_187_2 + shifted_state75_187_3);
      reservoir_sum_parallel[76] = (shifted_state76_1_0 + shifted_state76_1_1 + shifted_state76_1_2 + shifted_state76_1_5 + shifted_state76_1_6 + shifted_state76_1_7 + shifted_state76_2_2 + shifted_state76_2_4 + shifted_state76_14_5 + shifted_state76_33_4 + shifted_state76_35_0 + shifted_state76_35_1 + shifted_state76_35_3 + shifted_state76_35_4 + shifted_state76_35_6 + shifted_state76_35_7 + shifted_state76_42_0 + shifted_state76_42_2 + shifted_state76_42_4 + shifted_state76_42_5 + shifted_state76_42_6 + shifted_state76_42_7 + shifted_state76_71_2 + shifted_state76_71_4 + shifted_state76_71_5 + shifted_state76_71_6 + shifted_state76_71_7 + shifted_state76_73_0 + shifted_state76_73_4 + shifted_state76_74_0 + shifted_state76_74_3 + shifted_state76_95_0 + shifted_state76_95_4 + shifted_state76_95_6 + shifted_state76_95_7 + shifted_state76_99_1 + shifted_state76_99_2 + shifted_state76_99_3 + shifted_state76_99_6 + shifted_state76_99_7 + shifted_state76_121_1 + shifted_state76_121_2 + shifted_state76_121_3 + shifted_state76_121_5 + shifted_state76_129_4 + shifted_state76_129_6 + shifted_state76_129_7 + shifted_state76_154_0 + shifted_state76_154_2 + shifted_state76_154_3 + shifted_state76_154_4 + shifted_state76_154_6 + shifted_state76_154_7 + shifted_state76_159_0 + shifted_state76_159_1 + shifted_state76_159_3 + shifted_state76_159_5 + shifted_state76_164_0 + shifted_state76_164_2 + shifted_state76_164_3 + shifted_state76_164_6 + shifted_state76_164_7 + shifted_state76_172_0 + shifted_state76_172_5);
      reservoir_sum_parallel[77] = (shifted_state77_39_1 + shifted_state77_39_2 + shifted_state77_39_4 + shifted_state77_55_1 + shifted_state77_55_2 + shifted_state77_55_3 + shifted_state77_62_0 + shifted_state77_62_1 + shifted_state77_62_2 + shifted_state77_62_3 + shifted_state77_62_4 + shifted_state77_63_0 + shifted_state77_63_1 + shifted_state77_63_5 + shifted_state77_79_0 + shifted_state77_79_3 + shifted_state77_93_2 + shifted_state77_93_3 + shifted_state77_93_6 + shifted_state77_93_7 + shifted_state77_101_0 + shifted_state77_101_4 + shifted_state77_117_1 + shifted_state77_132_0 + shifted_state77_132_1 + shifted_state77_132_4 + shifted_state77_132_5 + shifted_state77_132_6 + shifted_state77_132_7 + shifted_state77_164_2 + shifted_state77_164_3 + shifted_state77_164_4 + shifted_state77_173_5 + shifted_state77_178_4 + shifted_state77_178_5 + shifted_state77_180_1 + shifted_state77_180_2 + shifted_state77_180_3 + shifted_state77_180_4 + shifted_state77_180_5);
      reservoir_sum_parallel[78] = (shifted_state78_21_1 + shifted_state78_21_2 + shifted_state78_21_6 + shifted_state78_30_1 + shifted_state78_30_3 + shifted_state78_45_0 + shifted_state78_45_1 + shifted_state78_45_5 + shifted_state78_45_6 + shifted_state78_45_7 + shifted_state78_48_0 + shifted_state78_52_0 + shifted_state78_52_2 + shifted_state78_52_3 + shifted_state78_52_5 + shifted_state78_52_6 + shifted_state78_52_7 + shifted_state78_83_0 + shifted_state78_83_2 + shifted_state78_83_3 + shifted_state78_83_4 + shifted_state78_83_5 + shifted_state78_83_6 + shifted_state78_83_7 + shifted_state78_90_1 + shifted_state78_90_2 + shifted_state78_90_6 + shifted_state78_90_7 + shifted_state78_103_0 + shifted_state78_103_1 + shifted_state78_112_1 + shifted_state78_112_4 + shifted_state78_112_6 + shifted_state78_112_7 + shifted_state78_122_1 + shifted_state78_125_2 + shifted_state78_125_3 + shifted_state78_128_2 + shifted_state78_128_4 + shifted_state78_128_5 + shifted_state78_128_6 + shifted_state78_128_7 + shifted_state78_133_0 + shifted_state78_133_3 + shifted_state78_133_4 + shifted_state78_133_6 + shifted_state78_133_7 + shifted_state78_142_3 + shifted_state78_162_1 + shifted_state78_162_2 + shifted_state78_162_3 + shifted_state78_162_4 + shifted_state78_162_5 + shifted_state78_162_6 + shifted_state78_162_7 + shifted_state78_171_4 + shifted_state78_171_5 + shifted_state78_181_0 + shifted_state78_181_4 + shifted_state78_181_5 + shifted_state78_192_0 + shifted_state78_192_1 + shifted_state78_192_3);
      reservoir_sum_parallel[79] = (shifted_state79_10_1 + shifted_state79_10_2 + shifted_state79_12_1 + shifted_state79_12_2 + shifted_state79_12_4 + shifted_state79_15_0 + shifted_state79_15_3 + shifted_state79_15_4 + shifted_state79_15_5 + shifted_state79_15_6 + shifted_state79_15_7 + shifted_state79_32_0 + shifted_state79_32_4 + shifted_state79_32_6 + shifted_state79_46_0 + shifted_state79_46_4 + shifted_state79_46_6 + shifted_state79_46_7 + shifted_state79_54_5 + shifted_state79_54_6 + shifted_state79_54_7 + shifted_state79_63_0 + shifted_state79_72_0 + shifted_state79_72_1 + shifted_state79_72_2 + shifted_state79_72_4 + shifted_state79_97_0 + shifted_state79_97_1 + shifted_state79_104_1 + shifted_state79_105_0 + shifted_state79_105_1 + shifted_state79_105_2 + shifted_state79_105_3 + shifted_state79_105_5 + shifted_state79_105_6 + shifted_state79_105_7 + shifted_state79_108_2 + shifted_state79_108_4 + shifted_state79_108_5 + shifted_state79_108_6 + shifted_state79_108_7 + shifted_state79_123_0 + shifted_state79_123_1 + shifted_state79_123_3 + shifted_state79_123_5 + shifted_state79_123_6 + shifted_state79_123_7 + shifted_state79_127_1 + shifted_state79_127_2 + shifted_state79_127_4 + shifted_state79_144_1 + shifted_state79_144_3 + shifted_state79_144_6 + shifted_state79_144_7 + shifted_state79_146_0 + shifted_state79_146_2 + shifted_state79_146_3 + shifted_state79_146_4 + shifted_state79_148_3 + shifted_state79_158_2 + shifted_state79_158_3 + shifted_state79_158_5 + shifted_state79_158_6 + shifted_state79_158_7 + shifted_state79_172_2 + shifted_state79_172_4 + shifted_state79_175_0 + shifted_state79_175_3 + shifted_state79_177_0 + shifted_state79_177_1 + shifted_state79_177_2 + shifted_state79_177_3 + shifted_state79_177_4 + shifted_state79_187_0 + shifted_state79_187_3 + shifted_state79_187_4 + shifted_state79_187_5 + shifted_state79_187_6 + shifted_state79_187_7 + shifted_state79_189_1 + shifted_state79_189_2 + shifted_state79_189_4 + shifted_state79_192_0 + shifted_state79_192_3 + shifted_state79_192_5);
      reservoir_sum_parallel[80] = (shifted_state80_24_1 + shifted_state80_25_1 + shifted_state80_25_2 + shifted_state80_25_4 + shifted_state80_25_5 + shifted_state80_25_6 + shifted_state80_25_7 + shifted_state80_37_0 + shifted_state80_37_1 + shifted_state80_37_2 + shifted_state80_37_5 + shifted_state80_37_6 + shifted_state80_37_7 + shifted_state80_40_0 + shifted_state80_40_1 + shifted_state80_40_4 + shifted_state80_40_6 + shifted_state80_40_7 + shifted_state80_48_0 + shifted_state80_48_1 + shifted_state80_48_2 + shifted_state80_48_3 + shifted_state80_52_1 + shifted_state80_52_2 + shifted_state80_52_3 + shifted_state80_52_4 + shifted_state80_52_6 + shifted_state80_52_7 + shifted_state80_57_1 + shifted_state80_57_2 + shifted_state80_57_3 + shifted_state80_57_4 + shifted_state80_57_5 + shifted_state80_57_6 + shifted_state80_57_7 + shifted_state80_67_0 + shifted_state80_67_3 + shifted_state80_67_4 + shifted_state80_67_5 + shifted_state80_67_6 + shifted_state80_67_7 + shifted_state80_77_0 + shifted_state80_77_1 + shifted_state80_77_2 + shifted_state80_77_3 + shifted_state80_77_4 + shifted_state80_86_0 + shifted_state80_86_4 + shifted_state80_92_0 + shifted_state80_92_1 + shifted_state80_92_3 + shifted_state80_94_0 + shifted_state80_94_1 + shifted_state80_94_2 + shifted_state80_94_3 + shifted_state80_115_2 + shifted_state80_115_3 + shifted_state80_115_5 + shifted_state80_126_0 + shifted_state80_126_1 + shifted_state80_126_5 + shifted_state80_153_0 + shifted_state80_153_4 + shifted_state80_153_5 + shifted_state80_153_6 + shifted_state80_153_7 + shifted_state80_158_0 + shifted_state80_158_1 + shifted_state80_158_4 + shifted_state80_158_5 + shifted_state80_158_6 + shifted_state80_158_7 + shifted_state80_163_0 + shifted_state80_163_1 + shifted_state80_163_3 + shifted_state80_163_4 + shifted_state80_163_5 + shifted_state80_163_6 + shifted_state80_163_7 + shifted_state80_164_1 + shifted_state80_166_0 + shifted_state80_166_1 + shifted_state80_166_3 + shifted_state80_166_4 + shifted_state80_168_1 + shifted_state80_168_2 + shifted_state80_168_3 + shifted_state80_168_4 + shifted_state80_175_1 + shifted_state80_175_3 + shifted_state80_177_2 + shifted_state80_177_4 + shifted_state80_189_0 + shifted_state80_191_1 + shifted_state80_191_3 + shifted_state80_191_5);
      reservoir_sum_parallel[81] = (shifted_state81_7_0 + shifted_state81_7_2 + shifted_state81_7_3 + shifted_state81_7_4 + shifted_state81_7_6 + shifted_state81_7_7 + shifted_state81_21_0 + shifted_state81_21_1 + shifted_state81_24_3 + shifted_state81_24_5 + shifted_state81_24_6 + shifted_state81_24_7 + shifted_state81_32_0 + shifted_state81_32_1 + shifted_state81_32_2 + shifted_state81_32_3 + shifted_state81_32_5 + shifted_state81_32_6 + shifted_state81_32_7 + shifted_state81_37_1 + shifted_state81_37_2 + shifted_state81_37_3 + shifted_state81_37_4 + shifted_state81_37_5 + shifted_state81_37_6 + shifted_state81_37_7 + shifted_state81_38_0 + shifted_state81_38_1 + shifted_state81_38_2 + shifted_state81_38_4 + shifted_state81_40_0 + shifted_state81_40_3 + shifted_state81_40_4 + shifted_state81_40_6 + shifted_state81_40_7 + shifted_state81_56_2 + shifted_state81_56_3 + shifted_state81_56_5 + shifted_state81_58_0 + shifted_state81_58_3 + shifted_state81_58_4 + shifted_state81_59_0 + shifted_state81_59_1 + shifted_state81_59_3 + shifted_state81_59_4 + shifted_state81_64_0 + shifted_state81_64_2 + shifted_state81_64_5 + shifted_state81_64_6 + shifted_state81_64_7 + shifted_state81_74_3 + shifted_state81_77_1 + shifted_state81_77_4 + shifted_state81_82_1 + shifted_state81_82_2 + shifted_state81_82_3 + shifted_state81_98_1 + shifted_state81_98_3 + shifted_state81_98_4 + shifted_state81_101_0 + shifted_state81_101_1 + shifted_state81_101_4 + shifted_state81_101_5 + shifted_state81_101_6 + shifted_state81_101_7 + shifted_state81_105_0 + shifted_state81_105_4 + shifted_state81_113_1 + shifted_state81_113_2 + shifted_state81_129_0 + shifted_state81_129_1 + shifted_state81_129_2 + shifted_state81_129_4 + shifted_state81_129_5 + shifted_state81_146_2 + shifted_state81_146_3 + shifted_state81_146_4 + shifted_state81_146_5 + shifted_state81_146_6 + shifted_state81_146_7 + shifted_state81_150_0 + shifted_state81_150_3 + shifted_state81_171_1 + shifted_state81_171_4 + shifted_state81_171_6 + shifted_state81_171_7 + shifted_state81_198_1 + shifted_state81_198_5);
      reservoir_sum_parallel[82] = (shifted_state82_7_3 + shifted_state82_7_4 + shifted_state82_8_0 + shifted_state82_8_1 + shifted_state82_12_0 + shifted_state82_12_1 + shifted_state82_12_3 + shifted_state82_15_2 + shifted_state82_15_3 + shifted_state82_29_1 + shifted_state82_38_0 + shifted_state82_38_1 + shifted_state82_38_3 + shifted_state82_41_0 + shifted_state82_41_1 + shifted_state82_41_2 + shifted_state82_41_5 + shifted_state82_60_0 + shifted_state82_60_5 + shifted_state82_60_6 + shifted_state82_60_7 + shifted_state82_72_3 + shifted_state82_72_4 + shifted_state82_72_5 + shifted_state82_72_6 + shifted_state82_72_7 + shifted_state82_74_1 + shifted_state82_74_2 + shifted_state82_74_5 + shifted_state82_74_6 + shifted_state82_74_7 + shifted_state82_91_2 + shifted_state82_91_3 + shifted_state82_91_4 + shifted_state82_91_5 + shifted_state82_91_6 + shifted_state82_91_7 + shifted_state82_104_0 + shifted_state82_104_1 + shifted_state82_104_3 + shifted_state82_104_5 + shifted_state82_104_6 + shifted_state82_104_7 + shifted_state82_129_0 + shifted_state82_129_2 + shifted_state82_129_3 + shifted_state82_136_0 + shifted_state82_136_2 + shifted_state82_136_3 + shifted_state82_136_4 + shifted_state82_146_0 + shifted_state82_146_1 + shifted_state82_146_4 + shifted_state82_146_5 + shifted_state82_146_6 + shifted_state82_146_7 + shifted_state82_149_0 + shifted_state82_149_1 + shifted_state82_149_2 + shifted_state82_149_3 + shifted_state82_149_4 + shifted_state82_149_5 + shifted_state82_149_7 + shifted_state82_154_2 + shifted_state82_154_3 + shifted_state82_154_4 + shifted_state82_154_5 + shifted_state82_154_6 + shifted_state82_154_7 + shifted_state82_167_0 + shifted_state82_167_1 + shifted_state82_167_2 + shifted_state82_167_3 + shifted_state82_167_4 + shifted_state82_167_6 + shifted_state82_167_7 + shifted_state82_170_0 + shifted_state82_170_1 + shifted_state82_170_3 + shifted_state82_170_4 + shifted_state82_170_5 + shifted_state82_170_7 + shifted_state82_188_0 + shifted_state82_188_1 + shifted_state82_188_3 + shifted_state82_188_4 + shifted_state82_188_6 + shifted_state82_188_7);
      reservoir_sum_parallel[83] = (shifted_state83_8_1 + shifted_state83_8_2 + shifted_state83_10_1 + shifted_state83_10_3 + shifted_state83_10_5 + shifted_state83_11_0 + shifted_state83_11_4 + shifted_state83_11_5 + shifted_state83_11_6 + shifted_state83_11_7 + shifted_state83_23_0 + shifted_state83_23_2 + shifted_state83_23_3 + shifted_state83_23_6 + shifted_state83_23_7 + shifted_state83_36_2 + shifted_state83_36_4 + shifted_state83_36_5 + shifted_state83_36_6 + shifted_state83_36_7 + shifted_state83_47_0 + shifted_state83_47_1 + shifted_state83_47_4 + shifted_state83_47_5 + shifted_state83_47_6 + shifted_state83_47_7 + shifted_state83_49_0 + shifted_state83_49_5 + shifted_state83_50_1 + shifted_state83_50_2 + shifted_state83_70_1 + shifted_state83_70_3 + shifted_state83_70_5 + shifted_state83_75_2 + shifted_state83_75_3 + shifted_state83_75_4 + shifted_state83_88_0 + shifted_state83_88_3 + shifted_state83_94_0 + shifted_state83_94_1 + shifted_state83_94_3 + shifted_state83_94_4 + shifted_state83_94_5 + shifted_state83_94_6 + shifted_state83_94_7 + shifted_state83_108_0 + shifted_state83_108_1 + shifted_state83_108_2 + shifted_state83_108_4 + shifted_state83_108_5 + shifted_state83_108_6 + shifted_state83_108_7 + shifted_state83_123_0 + shifted_state83_123_2 + shifted_state83_123_3 + shifted_state83_123_5 + shifted_state83_123_6 + shifted_state83_123_7 + shifted_state83_156_3 + shifted_state83_156_4);
      reservoir_sum_parallel[84] = (shifted_state84_5_2 + shifted_state84_5_3 + shifted_state84_22_0 + shifted_state84_22_4 + shifted_state84_28_1 + shifted_state84_28_4 + shifted_state84_70_1 + shifted_state84_70_3 + shifted_state84_70_4 + shifted_state84_70_5 + shifted_state84_70_7 + shifted_state84_74_0 + shifted_state84_74_1 + shifted_state84_74_5 + shifted_state84_78_0 + shifted_state84_79_3 + shifted_state84_79_4 + shifted_state84_79_5 + shifted_state84_79_6 + shifted_state84_79_7 + shifted_state84_80_1 + shifted_state84_80_2 + shifted_state84_80_3 + shifted_state84_80_4 + shifted_state84_80_5 + shifted_state84_80_6 + shifted_state84_80_7 + shifted_state84_91_0 + shifted_state84_91_4 + shifted_state84_91_5 + shifted_state84_91_6 + shifted_state84_91_7 + shifted_state84_109_1 + shifted_state84_109_2 + shifted_state84_109_3 + shifted_state84_109_4 + shifted_state84_109_5 + shifted_state84_109_6 + shifted_state84_109_7 + shifted_state84_114_0 + shifted_state84_114_3 + shifted_state84_122_0 + shifted_state84_122_1 + shifted_state84_122_3 + shifted_state84_122_5 + shifted_state84_122_6 + shifted_state84_122_7 + shifted_state84_136_5 + shifted_state84_136_6 + shifted_state84_136_7 + shifted_state84_157_3 + shifted_state84_157_5 + shifted_state84_157_6 + shifted_state84_157_7 + shifted_state84_167_0 + shifted_state84_167_1 + shifted_state84_167_2 + shifted_state84_194_1 + shifted_state84_194_5 + shifted_state84_194_6 + shifted_state84_194_7);
      reservoir_sum_parallel[85] = (shifted_state85_2_1 + shifted_state85_2_3 + shifted_state85_2_5 + shifted_state85_2_6 + shifted_state85_2_7 + shifted_state85_7_2 + shifted_state85_7_3 + shifted_state85_13_1 + shifted_state85_13_2 + shifted_state85_13_3 + shifted_state85_13_6 + shifted_state85_13_7 + shifted_state85_18_2 + shifted_state85_18_4 + shifted_state85_18_5 + shifted_state85_18_6 + shifted_state85_18_7 + shifted_state85_25_2 + shifted_state85_25_3 + shifted_state85_25_5 + shifted_state85_25_6 + shifted_state85_25_7 + shifted_state85_26_1 + shifted_state85_26_2 + shifted_state85_26_4 + shifted_state85_26_6 + shifted_state85_26_7 + shifted_state85_38_0 + shifted_state85_38_2 + shifted_state85_38_3 + shifted_state85_38_5 + shifted_state85_38_6 + shifted_state85_38_7 + shifted_state85_41_1 + shifted_state85_41_2 + shifted_state85_41_3 + shifted_state85_41_4 + shifted_state85_41_6 + shifted_state85_41_7 + shifted_state85_68_0 + shifted_state85_68_3 + shifted_state85_68_4 + shifted_state85_68_5 + shifted_state85_68_6 + shifted_state85_68_7 + shifted_state85_75_5 + shifted_state85_81_0 + shifted_state85_81_2 + shifted_state85_81_3 + shifted_state85_81_5 + shifted_state85_81_6 + shifted_state85_81_7 + shifted_state85_88_2 + shifted_state85_88_3 + shifted_state85_88_4 + shifted_state85_88_5 + shifted_state85_88_6 + shifted_state85_88_7 + shifted_state85_93_3 + shifted_state85_93_5 + shifted_state85_116_1 + shifted_state85_116_2 + shifted_state85_116_3 + shifted_state85_129_1 + shifted_state85_129_3 + shifted_state85_144_2 + shifted_state85_144_3 + shifted_state85_152_0 + shifted_state85_161_0 + shifted_state85_161_1 + shifted_state85_161_3 + shifted_state85_165_2 + shifted_state85_165_4 + shifted_state85_171_1 + shifted_state85_171_3 + shifted_state85_176_0 + shifted_state85_176_4 + shifted_state85_181_0 + shifted_state85_181_1 + shifted_state85_181_4 + shifted_state85_181_5 + shifted_state85_181_6 + shifted_state85_181_7 + shifted_state85_184_3 + shifted_state85_184_4 + shifted_state85_184_5 + shifted_state85_184_6 + shifted_state85_184_7 + shifted_state85_185_1 + shifted_state85_185_3 + shifted_state85_185_4 + shifted_state85_185_5 + shifted_state85_185_6 + shifted_state85_185_7 + shifted_state85_188_1 + shifted_state85_188_5 + shifted_state85_188_6 + shifted_state85_188_7 + shifted_state85_191_0 + shifted_state85_191_2 + shifted_state85_191_3 + shifted_state85_191_5 + shifted_state85_191_6 + shifted_state85_191_7 + shifted_state85_196_6);
      reservoir_sum_parallel[86] = (shifted_state86_3_0 + shifted_state86_3_3 + shifted_state86_3_5 + shifted_state86_3_6 + shifted_state86_3_7 + shifted_state86_9_0 + shifted_state86_9_1 + shifted_state86_9_2 + shifted_state86_9_3 + shifted_state86_9_5 + shifted_state86_9_6 + shifted_state86_9_7 + shifted_state86_18_3 + shifted_state86_40_4 + shifted_state86_40_5 + shifted_state86_40_6 + shifted_state86_40_7 + shifted_state86_50_0 + shifted_state86_50_1 + shifted_state86_50_2 + shifted_state86_50_5 + shifted_state86_54_1 + shifted_state86_54_2 + shifted_state86_55_0 + shifted_state86_55_1 + shifted_state86_55_3 + shifted_state86_55_4 + shifted_state86_55_6 + shifted_state86_55_7 + shifted_state86_63_0 + shifted_state86_63_2 + shifted_state86_63_5 + shifted_state86_63_6 + shifted_state86_63_7 + shifted_state86_76_0 + shifted_state86_76_2 + shifted_state86_76_4 + shifted_state86_76_6 + shifted_state86_76_7 + shifted_state86_80_0 + shifted_state86_80_1 + shifted_state86_80_2 + shifted_state86_80_3 + shifted_state86_80_5 + shifted_state86_80_6 + shifted_state86_80_7 + shifted_state86_88_1 + shifted_state86_88_2 + shifted_state86_88_3 + shifted_state86_88_4 + shifted_state86_88_6 + shifted_state86_88_7 + shifted_state86_93_0 + shifted_state86_93_3 + shifted_state86_93_5 + shifted_state86_93_6 + shifted_state86_93_7 + shifted_state86_105_1 + shifted_state86_105_4 + shifted_state86_105_5 + shifted_state86_105_6 + shifted_state86_105_7 + shifted_state86_109_0 + shifted_state86_109_2 + shifted_state86_109_3 + shifted_state86_118_1 + shifted_state86_118_2 + shifted_state86_118_3 + shifted_state86_118_4 + shifted_state86_118_5 + shifted_state86_118_7 + shifted_state86_131_0 + shifted_state86_131_3 + shifted_state86_131_5 + shifted_state86_131_6 + shifted_state86_131_7 + shifted_state86_137_2 + shifted_state86_137_5 + shifted_state86_139_1 + shifted_state86_139_2 + shifted_state86_139_5 + shifted_state86_139_6 + shifted_state86_139_7 + shifted_state86_141_1 + shifted_state86_141_4 + shifted_state86_141_5 + shifted_state86_141_6 + shifted_state86_141_7 + shifted_state86_153_0 + shifted_state86_153_1 + shifted_state86_153_4 + shifted_state86_164_0 + shifted_state86_164_1 + shifted_state86_164_6 + shifted_state86_167_2 + shifted_state86_167_5 + shifted_state86_167_7 + shifted_state86_168_0 + shifted_state86_168_1 + shifted_state86_168_3 + shifted_state86_169_1 + shifted_state86_169_2 + shifted_state86_169_3 + shifted_state86_169_5 + shifted_state86_169_6 + shifted_state86_169_7 + shifted_state86_171_2 + shifted_state86_180_1 + shifted_state86_180_2 + shifted_state86_180_3 + shifted_state86_180_5 + shifted_state86_180_6 + shifted_state86_180_7 + shifted_state86_188_2 + shifted_state86_188_3 + shifted_state86_188_4 + shifted_state86_195_1 + shifted_state86_195_2 + shifted_state86_195_4 + shifted_state86_195_5 + shifted_state86_198_0 + shifted_state86_198_1 + shifted_state86_198_4 + shifted_state86_198_5 + shifted_state86_198_7 + shifted_state86_199_0 + shifted_state86_199_1 + shifted_state86_199_4);
      reservoir_sum_parallel[87] = (shifted_state87_0_4 + shifted_state87_7_2 + shifted_state87_7_4 + shifted_state87_7_5 + shifted_state87_7_6 + shifted_state87_7_7 + shifted_state87_12_1 + shifted_state87_12_2 + shifted_state87_12_6 + shifted_state87_23_0 + shifted_state87_23_1 + shifted_state87_23_2 + shifted_state87_26_1 + shifted_state87_26_2 + shifted_state87_26_4 + shifted_state87_26_5 + shifted_state87_26_6 + shifted_state87_26_7 + shifted_state87_38_4 + shifted_state87_40_0 + shifted_state87_40_1 + shifted_state87_40_2 + shifted_state87_40_3 + shifted_state87_48_0 + shifted_state87_48_1 + shifted_state87_48_2 + shifted_state87_48_3 + shifted_state87_48_5 + shifted_state87_49_0 + shifted_state87_49_2 + shifted_state87_49_5 + shifted_state87_50_0 + shifted_state87_60_0 + shifted_state87_60_1 + shifted_state87_60_3 + shifted_state87_60_4 + shifted_state87_67_0 + shifted_state87_67_1 + shifted_state87_67_2 + shifted_state87_67_3 + shifted_state87_67_5 + shifted_state87_74_2 + shifted_state87_74_5 + shifted_state87_74_6 + shifted_state87_74_7 + shifted_state87_93_0 + shifted_state87_93_1 + shifted_state87_93_2 + shifted_state87_93_6 + shifted_state87_101_2 + shifted_state87_101_4 + shifted_state87_101_6 + shifted_state87_101_7 + shifted_state87_103_1 + shifted_state87_103_2 + shifted_state87_103_5 + shifted_state87_103_6 + shifted_state87_103_7 + shifted_state87_108_0 + shifted_state87_108_3 + shifted_state87_111_2 + shifted_state87_111_3 + shifted_state87_111_5 + shifted_state87_113_1 + shifted_state87_113_2 + shifted_state87_121_4 + shifted_state87_121_5 + shifted_state87_121_6 + shifted_state87_121_7 + shifted_state87_131_0 + shifted_state87_131_1 + shifted_state87_131_3 + shifted_state87_131_4 + shifted_state87_131_5 + shifted_state87_131_6 + shifted_state87_131_7 + shifted_state87_141_0 + shifted_state87_141_6 + shifted_state87_141_7 + shifted_state87_152_0 + shifted_state87_152_1 + shifted_state87_152_2 + shifted_state87_152_4 + shifted_state87_152_5 + shifted_state87_153_2 + shifted_state87_153_4 + shifted_state87_155_3 + shifted_state87_155_4 + shifted_state87_155_5 + shifted_state87_157_5 + shifted_state87_191_0 + shifted_state87_191_1 + shifted_state87_191_2 + shifted_state87_191_4);
      reservoir_sum_parallel[88] = (shifted_state88_1_0 + shifted_state88_1_1 + shifted_state88_1_2 + shifted_state88_1_3 + shifted_state88_1_4 + shifted_state88_1_5 + shifted_state88_1_6 + shifted_state88_1_7 + shifted_state88_5_0 + shifted_state88_5_3 + shifted_state88_8_0 + shifted_state88_8_2 + shifted_state88_8_4 + shifted_state88_10_1 + shifted_state88_10_3 + shifted_state88_10_4 + shifted_state88_10_6 + shifted_state88_10_7 + shifted_state88_13_0 + shifted_state88_13_2 + shifted_state88_13_4 + shifted_state88_13_5 + shifted_state88_13_6 + shifted_state88_13_7 + shifted_state88_45_0 + shifted_state88_45_1 + shifted_state88_45_2 + shifted_state88_45_5 + shifted_state88_74_3 + shifted_state88_74_4 + shifted_state88_92_1 + shifted_state88_92_3 + shifted_state88_92_4 + shifted_state88_103_1 + shifted_state88_103_3 + shifted_state88_103_5 + shifted_state88_103_6 + shifted_state88_103_7 + shifted_state88_123_2 + shifted_state88_123_5 + shifted_state88_123_6 + shifted_state88_123_7 + shifted_state88_130_0 + shifted_state88_130_3 + shifted_state88_130_4 + shifted_state88_154_1 + shifted_state88_154_2 + shifted_state88_154_4 + shifted_state88_154_5 + shifted_state88_154_6 + shifted_state88_154_7 + shifted_state88_162_1 + shifted_state88_162_4 + shifted_state88_163_2 + shifted_state88_167_0 + shifted_state88_167_5 + shifted_state88_183_0 + shifted_state88_183_2 + shifted_state88_183_3 + shifted_state88_193_0 + shifted_state88_193_2 + shifted_state88_193_4 + shifted_state88_197_3 + shifted_state88_197_4 + shifted_state88_197_5 + shifted_state88_197_6 + shifted_state88_197_7);
      reservoir_sum_parallel[89] = (shifted_state89_6_0 + shifted_state89_6_2 + shifted_state89_6_4 + shifted_state89_13_0 + shifted_state89_13_2 + shifted_state89_16_0 + shifted_state89_16_1 + shifted_state89_16_5 + shifted_state89_16_6 + shifted_state89_16_7 + shifted_state89_19_0 + shifted_state89_19_2 + shifted_state89_19_3 + shifted_state89_19_4 + shifted_state89_28_0 + shifted_state89_28_2 + shifted_state89_28_3 + shifted_state89_50_0 + shifted_state89_50_2 + shifted_state89_50_4 + shifted_state89_58_1 + shifted_state89_58_4 + shifted_state89_58_6 + shifted_state89_58_7 + shifted_state89_64_1 + shifted_state89_64_2 + shifted_state89_71_0 + shifted_state89_71_2 + shifted_state89_71_3 + shifted_state89_71_4 + shifted_state89_71_5 + shifted_state89_71_6 + shifted_state89_71_7 + shifted_state89_74_0 + shifted_state89_74_4 + shifted_state89_78_0 + shifted_state89_78_5 + shifted_state89_79_0 + shifted_state89_79_2 + shifted_state89_79_4 + shifted_state89_79_5 + shifted_state89_79_6 + shifted_state89_79_7 + shifted_state89_80_3 + shifted_state89_93_3 + shifted_state89_93_5 + shifted_state89_93_6 + shifted_state89_93_7 + shifted_state89_122_0 + shifted_state89_122_1 + shifted_state89_122_2 + shifted_state89_122_3 + shifted_state89_122_4 + shifted_state89_122_6 + shifted_state89_122_7 + shifted_state89_126_0 + shifted_state89_126_2 + shifted_state89_134_0 + shifted_state89_134_1 + shifted_state89_134_3 + shifted_state89_134_4 + shifted_state89_142_2 + shifted_state89_142_3 + shifted_state89_144_0 + shifted_state89_144_1 + shifted_state89_144_5 + shifted_state89_153_1 + shifted_state89_153_3 + shifted_state89_153_5 + shifted_state89_153_6 + shifted_state89_153_7 + shifted_state89_156_2 + shifted_state89_156_3 + shifted_state89_156_5 + shifted_state89_176_1 + shifted_state89_176_2 + shifted_state89_176_3 + shifted_state89_177_3 + shifted_state89_177_5 + shifted_state89_177_6 + shifted_state89_177_7 + shifted_state89_181_1 + shifted_state89_181_2 + shifted_state89_181_4 + shifted_state89_182_3 + shifted_state89_182_4 + shifted_state89_182_5 + shifted_state89_182_6 + shifted_state89_182_7 + shifted_state89_188_1 + shifted_state89_188_3 + shifted_state89_188_5 + shifted_state89_188_6 + shifted_state89_188_7 + shifted_state89_189_1 + shifted_state89_189_2 + shifted_state89_189_3 + shifted_state89_189_5 + shifted_state89_189_6 + shifted_state89_189_7);
      reservoir_sum_parallel[90] = (shifted_state90_4_0 + shifted_state90_4_1 + shifted_state90_4_3 + shifted_state90_4_4 + shifted_state90_4_6 + shifted_state90_4_7 + shifted_state90_6_1 + shifted_state90_6_2 + shifted_state90_6_3 + shifted_state90_6_4 + shifted_state90_6_6 + shifted_state90_6_7 + shifted_state90_13_2 + shifted_state90_13_6 + shifted_state90_19_1 + shifted_state90_19_2 + shifted_state90_19_4 + shifted_state90_19_5 + shifted_state90_19_6 + shifted_state90_19_7 + shifted_state90_33_0 + shifted_state90_33_2 + shifted_state90_33_5 + shifted_state90_33_6 + shifted_state90_33_7 + shifted_state90_69_0 + shifted_state90_69_1 + shifted_state90_69_2 + shifted_state90_69_3 + shifted_state90_69_4 + shifted_state90_69_6 + shifted_state90_69_7 + shifted_state90_100_1 + shifted_state90_100_2 + shifted_state90_114_0 + shifted_state90_114_1 + shifted_state90_114_3 + shifted_state90_114_4 + shifted_state90_117_4 + shifted_state90_117_5 + shifted_state90_122_0 + shifted_state90_122_1 + shifted_state90_122_2 + shifted_state90_122_5 + shifted_state90_130_0 + shifted_state90_138_1 + shifted_state90_138_2 + shifted_state90_138_3 + shifted_state90_138_4 + shifted_state90_152_2 + shifted_state90_152_3 + shifted_state90_155_1 + shifted_state90_155_5 + shifted_state90_167_4 + shifted_state90_167_5 + shifted_state90_167_6 + shifted_state90_167_7 + shifted_state90_178_0 + shifted_state90_178_2 + shifted_state90_178_3);
      reservoir_sum_parallel[91] = (shifted_state91_3_0 + shifted_state91_3_1 + shifted_state91_3_3 + shifted_state91_20_4 + shifted_state91_20_5 + shifted_state91_20_6 + shifted_state91_20_7 + shifted_state91_29_0 + shifted_state91_29_2 + shifted_state91_29_6 + shifted_state91_29_7 + shifted_state91_47_1 + shifted_state91_47_3 + shifted_state91_47_6 + shifted_state91_56_0 + shifted_state91_56_2 + shifted_state91_56_3 + shifted_state91_56_6 + shifted_state91_56_7 + shifted_state91_64_0 + shifted_state91_64_3 + shifted_state91_64_4 + shifted_state91_64_6 + shifted_state91_64_7 + shifted_state91_73_3 + shifted_state91_73_5 + shifted_state91_73_6 + shifted_state91_73_7 + shifted_state91_87_0 + shifted_state91_87_1 + shifted_state91_87_3 + shifted_state91_87_4 + shifted_state91_87_5 + shifted_state91_87_6 + shifted_state91_87_7 + shifted_state91_93_0 + shifted_state91_93_1 + shifted_state91_93_3 + shifted_state91_96_0 + shifted_state91_96_1 + shifted_state91_96_2 + shifted_state91_96_4 + shifted_state91_96_5 + shifted_state91_96_6 + shifted_state91_96_7 + shifted_state91_103_1 + shifted_state91_103_2 + shifted_state91_103_3 + shifted_state91_103_5 + shifted_state91_103_6 + shifted_state91_103_7 + shifted_state91_104_3 + shifted_state91_104_4 + shifted_state91_104_5 + shifted_state91_104_6 + shifted_state91_104_7 + shifted_state91_109_2 + shifted_state91_118_0 + shifted_state91_142_1 + shifted_state91_142_3 + shifted_state91_142_4 + shifted_state91_142_6 + shifted_state91_142_7 + shifted_state91_150_0 + shifted_state91_150_1 + shifted_state91_150_4 + shifted_state91_150_6 + shifted_state91_150_7 + shifted_state91_166_1 + shifted_state91_174_0 + shifted_state91_174_1 + shifted_state91_174_3 + shifted_state91_183_1 + shifted_state91_183_5 + shifted_state91_184_0 + shifted_state91_184_2 + shifted_state91_189_1 + shifted_state91_189_3 + shifted_state91_189_4 + shifted_state91_189_5 + shifted_state91_194_0 + shifted_state91_194_1 + shifted_state91_194_2 + shifted_state91_194_3 + shifted_state91_194_5 + shifted_state91_194_6 + shifted_state91_194_7);
      reservoir_sum_parallel[92] = (shifted_state92_16_0 + shifted_state92_16_2 + shifted_state92_18_2 + shifted_state92_18_3 + shifted_state92_18_4 + shifted_state92_21_2 + shifted_state92_39_0 + shifted_state92_39_1 + shifted_state92_39_2 + shifted_state92_39_3 + shifted_state92_39_4 + shifted_state92_71_0 + shifted_state92_74_4 + shifted_state92_74_5 + shifted_state92_74_6 + shifted_state92_74_7 + shifted_state92_84_0 + shifted_state92_84_1 + shifted_state92_84_2 + shifted_state92_84_3 + shifted_state92_84_4 + shifted_state92_84_5 + shifted_state92_84_6 + shifted_state92_84_7 + shifted_state92_93_1 + shifted_state92_100_0 + shifted_state92_100_2 + shifted_state92_100_5 + shifted_state92_103_1 + shifted_state92_103_2 + shifted_state92_105_3 + shifted_state92_105_5 + shifted_state92_119_0 + shifted_state92_119_1 + shifted_state92_119_3 + shifted_state92_119_4 + shifted_state92_119_6 + shifted_state92_119_7 + shifted_state92_121_3 + shifted_state92_121_4 + shifted_state92_121_5 + shifted_state92_126_1 + shifted_state92_126_2 + shifted_state92_126_4 + shifted_state92_126_6 + shifted_state92_126_7 + shifted_state92_137_0 + shifted_state92_137_1 + shifted_state92_137_2 + shifted_state92_137_3 + shifted_state92_137_4 + shifted_state92_137_5 + shifted_state92_137_6 + shifted_state92_137_7 + shifted_state92_141_3 + shifted_state92_145_2 + shifted_state92_155_0 + shifted_state92_155_1 + shifted_state92_155_2 + shifted_state92_173_0 + shifted_state92_173_1 + shifted_state92_173_2 + shifted_state92_173_4 + shifted_state92_173_6 + shifted_state92_173_7 + shifted_state92_193_1 + shifted_state92_193_2 + shifted_state92_193_4 + shifted_state92_193_5);
      reservoir_sum_parallel[93] = (shifted_state93_9_0 + shifted_state93_9_1 + shifted_state93_9_3 + shifted_state93_9_4 + shifted_state93_9_5 + shifted_state93_9_6 + shifted_state93_9_7 + shifted_state93_27_1 + shifted_state93_27_2 + shifted_state93_27_3 + shifted_state93_27_6 + shifted_state93_27_7 + shifted_state93_44_1 + shifted_state93_44_2 + shifted_state93_44_4 + shifted_state93_44_5 + shifted_state93_44_6 + shifted_state93_44_7 + shifted_state93_61_0 + shifted_state93_61_3 + shifted_state93_61_4 + shifted_state93_61_5 + shifted_state93_61_6 + shifted_state93_61_7 + shifted_state93_80_2 + shifted_state93_80_3 + shifted_state93_80_4 + shifted_state93_83_0 + shifted_state93_83_1 + shifted_state93_83_2 + shifted_state93_83_3 + shifted_state93_83_4 + shifted_state93_83_5 + shifted_state93_83_6 + shifted_state93_83_7 + shifted_state93_100_0 + shifted_state93_100_1 + shifted_state93_100_2 + shifted_state93_100_3 + shifted_state93_100_4 + shifted_state93_100_6 + shifted_state93_104_0 + shifted_state93_104_4 + shifted_state93_104_5 + shifted_state93_104_6 + shifted_state93_104_7 + shifted_state93_107_0 + shifted_state93_107_1 + shifted_state93_107_2 + shifted_state93_107_4 + shifted_state93_107_5 + shifted_state93_107_6 + shifted_state93_107_7 + shifted_state93_112_0 + shifted_state93_112_1 + shifted_state93_112_3 + shifted_state93_123_1 + shifted_state93_123_5 + shifted_state93_123_6 + shifted_state93_123_7 + shifted_state93_126_1 + shifted_state93_126_5 + shifted_state93_126_6 + shifted_state93_126_7 + shifted_state93_143_1 + shifted_state93_143_2 + shifted_state93_143_5 + shifted_state93_143_6 + shifted_state93_143_7 + shifted_state93_149_0 + shifted_state93_149_2 + shifted_state93_149_3 + shifted_state93_149_5 + shifted_state93_150_1 + shifted_state93_150_2 + shifted_state93_150_3 + shifted_state93_150_4 + shifted_state93_150_5 + shifted_state93_150_6 + shifted_state93_150_7 + shifted_state93_151_0 + shifted_state93_151_2 + shifted_state93_151_4 + shifted_state93_170_0 + shifted_state93_170_1 + shifted_state93_170_2 + shifted_state93_170_3 + shifted_state93_170_5 + shifted_state93_170_6 + shifted_state93_170_7 + shifted_state93_180_0 + shifted_state93_180_4 + shifted_state93_180_5 + shifted_state93_180_6 + shifted_state93_180_7 + shifted_state93_181_0 + shifted_state93_181_2 + shifted_state93_181_5 + shifted_state93_181_6 + shifted_state93_181_7 + shifted_state93_185_1 + shifted_state93_185_2);
      reservoir_sum_parallel[94] = (shifted_state94_2_0 + shifted_state94_2_2 + shifted_state94_2_3 + shifted_state94_2_4 + shifted_state94_2_5 + shifted_state94_2_6 + shifted_state94_2_7 + shifted_state94_11_2 + shifted_state94_11_3 + shifted_state94_11_4 + shifted_state94_18_0 + shifted_state94_18_4 + shifted_state94_18_5 + shifted_state94_26_0 + shifted_state94_26_1 + shifted_state94_26_4 + shifted_state94_26_5 + shifted_state94_26_6 + shifted_state94_26_7 + shifted_state94_28_0 + shifted_state94_28_1 + shifted_state94_28_4 + shifted_state94_28_6 + shifted_state94_28_7 + shifted_state94_37_1 + shifted_state94_37_3 + shifted_state94_37_5 + shifted_state94_50_1 + shifted_state94_50_2 + shifted_state94_50_3 + shifted_state94_50_5 + shifted_state94_50_6 + shifted_state94_50_7 + shifted_state94_57_5 + shifted_state94_63_1 + shifted_state94_63_2 + shifted_state94_63_3 + shifted_state94_63_5 + shifted_state94_63_6 + shifted_state94_63_7 + shifted_state94_71_2 + shifted_state94_71_5 + shifted_state94_84_5 + shifted_state94_91_0 + shifted_state94_91_4 + shifted_state94_96_1 + shifted_state94_96_2 + shifted_state94_96_4 + shifted_state94_102_1 + shifted_state94_102_2 + shifted_state94_102_5 + shifted_state94_102_6 + shifted_state94_102_7 + shifted_state94_121_0 + shifted_state94_121_2 + shifted_state94_121_5 + shifted_state94_121_6 + shifted_state94_127_1 + shifted_state94_127_5 + shifted_state94_127_6 + shifted_state94_127_7 + shifted_state94_179_4 + shifted_state94_179_5 + shifted_state94_179_6 + shifted_state94_179_7 + shifted_state94_182_3 + shifted_state94_182_4 + shifted_state94_187_0 + shifted_state94_187_2 + shifted_state94_187_3 + shifted_state94_187_4 + shifted_state94_187_6 + shifted_state94_187_7 + shifted_state94_192_1 + shifted_state94_192_5 + shifted_state94_194_4 + shifted_state94_194_5 + shifted_state94_194_6 + shifted_state94_194_7);
      reservoir_sum_parallel[95] = (shifted_state95_0_0 + shifted_state95_0_1 + shifted_state95_0_2 + shifted_state95_0_4 + shifted_state95_0_6 + shifted_state95_0_7 + shifted_state95_30_2 + shifted_state95_30_3 + shifted_state95_30_5 + shifted_state95_30_6 + shifted_state95_30_7 + shifted_state95_39_2 + shifted_state95_39_4 + shifted_state95_39_5 + shifted_state95_39_6 + shifted_state95_39_7 + shifted_state95_61_2 + shifted_state95_61_3 + shifted_state95_73_0 + shifted_state95_73_2 + shifted_state95_73_4 + shifted_state95_78_0 + shifted_state95_78_2 + shifted_state95_78_4 + shifted_state95_98_2 + shifted_state95_98_4 + shifted_state95_98_5 + shifted_state95_98_6 + shifted_state95_98_7 + shifted_state95_107_0 + shifted_state95_107_4 + shifted_state95_111_1 + shifted_state95_111_3 + shifted_state95_111_6 + shifted_state95_111_7 + shifted_state95_117_0 + shifted_state95_117_1 + shifted_state95_117_2 + shifted_state95_117_3 + shifted_state95_147_0 + shifted_state95_147_1 + shifted_state95_147_2 + shifted_state95_147_3 + shifted_state95_147_4 + shifted_state95_149_0 + shifted_state95_149_4 + shifted_state95_149_5 + shifted_state95_159_0 + shifted_state95_159_3 + shifted_state95_159_4 + shifted_state95_161_1 + shifted_state95_161_2 + shifted_state95_161_3 + shifted_state95_161_4 + shifted_state95_161_5 + shifted_state95_161_6 + shifted_state95_161_7 + shifted_state95_166_0 + shifted_state95_166_2 + shifted_state95_166_3 + shifted_state95_166_4 + shifted_state95_166_5 + shifted_state95_166_6 + shifted_state95_166_7 + shifted_state95_171_0 + shifted_state95_171_1 + shifted_state95_172_0 + shifted_state95_176_1 + shifted_state95_176_3 + shifted_state95_176_5 + shifted_state95_176_6 + shifted_state95_176_7 + shifted_state95_179_0 + shifted_state95_179_1 + shifted_state95_179_3 + shifted_state95_179_5 + shifted_state95_179_6 + shifted_state95_179_7);
      reservoir_sum_parallel[96] = (shifted_state96_3_0 + shifted_state96_3_1 + shifted_state96_3_2 + shifted_state96_3_4 + shifted_state96_3_5 + shifted_state96_19_3 + shifted_state96_22_0 + shifted_state96_22_2 + shifted_state96_22_3 + shifted_state96_22_4 + shifted_state96_22_5 + shifted_state96_22_6 + shifted_state96_22_7 + shifted_state96_28_1 + shifted_state96_28_2 + shifted_state96_28_3 + shifted_state96_28_5 + shifted_state96_28_6 + shifted_state96_28_7 + shifted_state96_42_1 + shifted_state96_42_4 + shifted_state96_42_5 + shifted_state96_48_1 + shifted_state96_48_3 + shifted_state96_48_5 + shifted_state96_48_6 + shifted_state96_48_7 + shifted_state96_49_0 + shifted_state96_49_1 + shifted_state96_49_4 + shifted_state96_49_5 + shifted_state96_49_6 + shifted_state96_49_7 + shifted_state96_52_2 + shifted_state96_52_3 + shifted_state96_52_5 + shifted_state96_63_0 + shifted_state96_63_1 + shifted_state96_63_2 + shifted_state96_63_3 + shifted_state96_63_6 + shifted_state96_63_7 + shifted_state96_80_0 + shifted_state96_80_1 + shifted_state96_80_3 + shifted_state96_80_5 + shifted_state96_80_6 + shifted_state96_80_7 + shifted_state96_85_1 + shifted_state96_85_4 + shifted_state96_106_0 + shifted_state96_106_1 + shifted_state96_106_3 + shifted_state96_106_5 + shifted_state96_106_6 + shifted_state96_106_7 + shifted_state96_129_0 + shifted_state96_129_1 + shifted_state96_129_2 + shifted_state96_129_4 + shifted_state96_129_5 + shifted_state96_129_6 + shifted_state96_129_7 + shifted_state96_133_1 + shifted_state96_133_3 + shifted_state96_139_0 + shifted_state96_139_1 + shifted_state96_139_3 + shifted_state96_139_4 + shifted_state96_139_6 + shifted_state96_139_7 + shifted_state96_173_0 + shifted_state96_173_2 + shifted_state96_173_3 + shifted_state96_173_4 + shifted_state96_173_5 + shifted_state96_173_6 + shifted_state96_173_7);
      reservoir_sum_parallel[97] = (shifted_state97_4_1 + shifted_state97_4_2 + shifted_state97_6_0 + shifted_state97_6_1 + shifted_state97_6_2 + shifted_state97_6_5 + shifted_state97_6_6 + shifted_state97_6_7 + shifted_state97_31_1 + shifted_state97_31_2 + shifted_state97_31_5 + shifted_state97_31_6 + shifted_state97_31_7 + shifted_state97_34_1 + shifted_state97_34_4 + shifted_state97_46_0 + shifted_state97_46_4 + shifted_state97_46_6 + shifted_state97_46_7 + shifted_state97_63_1 + shifted_state97_63_3 + shifted_state97_63_6 + shifted_state97_63_7 + shifted_state97_71_1 + shifted_state97_71_4 + shifted_state97_71_5 + shifted_state97_71_6 + shifted_state97_71_7 + shifted_state97_89_0 + shifted_state97_89_1 + shifted_state97_89_3 + shifted_state97_135_0 + shifted_state97_135_3 + shifted_state97_135_6 + shifted_state97_135_7 + shifted_state97_141_0 + shifted_state97_164_0 + shifted_state97_164_1 + shifted_state97_164_2 + shifted_state97_164_4 + shifted_state97_164_5 + shifted_state97_166_0 + shifted_state97_166_5 + shifted_state97_167_0 + shifted_state97_167_1 + shifted_state97_167_2 + shifted_state97_167_5 + shifted_state97_167_6 + shifted_state97_167_7 + shifted_state97_168_0 + shifted_state97_168_1 + shifted_state97_168_3 + shifted_state97_168_4 + shifted_state97_168_6 + shifted_state97_168_7 + shifted_state97_170_4 + shifted_state97_195_2);
      reservoir_sum_parallel[98] = (shifted_state98_7_1 + shifted_state98_7_4 + shifted_state98_7_6 + shifted_state98_7_7 + shifted_state98_10_2 + shifted_state98_10_3 + shifted_state98_10_4 + shifted_state98_35_0 + shifted_state98_38_1 + shifted_state98_38_3 + shifted_state98_43_1 + shifted_state98_43_2 + shifted_state98_43_3 + shifted_state98_43_5 + shifted_state98_50_0 + shifted_state98_50_1 + shifted_state98_54_0 + shifted_state98_54_6 + shifted_state98_68_3 + shifted_state98_68_4 + shifted_state98_72_1 + shifted_state98_72_2 + shifted_state98_72_3 + shifted_state98_72_4 + shifted_state98_72_5 + shifted_state98_72_6 + shifted_state98_72_7 + shifted_state98_75_0 + shifted_state98_75_1 + shifted_state98_75_2 + shifted_state98_77_1 + shifted_state98_77_2 + shifted_state98_77_6 + shifted_state98_77_7 + shifted_state98_86_3 + shifted_state98_86_5 + shifted_state98_91_2 + shifted_state98_91_4 + shifted_state98_91_5 + shifted_state98_91_6 + shifted_state98_91_7 + shifted_state98_97_0 + shifted_state98_97_1 + shifted_state98_97_2 + shifted_state98_97_3 + shifted_state98_97_5 + shifted_state98_97_6 + shifted_state98_97_7 + shifted_state98_99_3 + shifted_state98_99_5 + shifted_state98_102_0 + shifted_state98_102_5 + shifted_state98_108_0 + shifted_state98_108_1 + shifted_state98_108_2 + shifted_state98_108_3 + shifted_state98_108_6 + shifted_state98_108_7 + shifted_state98_115_0 + shifted_state98_115_1 + shifted_state98_115_3 + shifted_state98_115_4 + shifted_state98_115_5 + shifted_state98_115_6 + shifted_state98_115_7 + shifted_state98_118_0 + shifted_state98_118_1 + shifted_state98_119_0 + shifted_state98_119_2 + shifted_state98_119_4 + shifted_state98_119_5 + shifted_state98_119_6 + shifted_state98_119_7 + shifted_state98_133_0 + shifted_state98_133_1 + shifted_state98_133_5 + shifted_state98_139_2 + shifted_state98_139_3 + shifted_state98_139_5 + shifted_state98_139_6 + shifted_state98_139_7 + shifted_state98_140_5 + shifted_state98_140_6 + shifted_state98_140_7 + shifted_state98_170_0 + shifted_state98_170_2 + shifted_state98_170_4 + shifted_state98_177_3 + shifted_state98_192_0 + shifted_state98_192_4 + shifted_state98_196_0 + shifted_state98_196_1 + shifted_state98_196_3 + shifted_state98_196_4 + shifted_state98_198_0 + shifted_state98_198_2 + shifted_state98_198_3 + shifted_state98_198_4 + shifted_state98_198_5);
      reservoir_sum_parallel[99] = (shifted_state99_0_0 + shifted_state99_0_1 + shifted_state99_0_2 + shifted_state99_0_3 + shifted_state99_0_4 + shifted_state99_0_6 + shifted_state99_0_7 + shifted_state99_2_1 + shifted_state99_2_2 + shifted_state99_2_3 + shifted_state99_2_4 + shifted_state99_2_5 + shifted_state99_2_6 + shifted_state99_2_7 + shifted_state99_26_0 + shifted_state99_26_1 + shifted_state99_26_5 + shifted_state99_26_6 + shifted_state99_26_7 + shifted_state99_31_0 + shifted_state99_31_2 + shifted_state99_31_4 + shifted_state99_31_5 + shifted_state99_31_6 + shifted_state99_31_7 + shifted_state99_50_1 + shifted_state99_50_3 + shifted_state99_50_6 + shifted_state99_50_7 + shifted_state99_56_2 + shifted_state99_56_4 + shifted_state99_56_5 + shifted_state99_56_6 + shifted_state99_56_7 + shifted_state99_59_0 + shifted_state99_59_1 + shifted_state99_59_4 + shifted_state99_76_0 + shifted_state99_76_4 + shifted_state99_76_5 + shifted_state99_76_6 + shifted_state99_76_7 + shifted_state99_77_0 + shifted_state99_77_3 + shifted_state99_77_4 + shifted_state99_77_5 + shifted_state99_77_7 + shifted_state99_84_0 + shifted_state99_86_0 + shifted_state99_86_1 + shifted_state99_90_3 + shifted_state99_90_4 + shifted_state99_90_6 + shifted_state99_90_7 + shifted_state99_96_0 + shifted_state99_96_2 + shifted_state99_96_3 + shifted_state99_96_5 + shifted_state99_96_6 + shifted_state99_96_7 + shifted_state99_101_0 + shifted_state99_101_1 + shifted_state99_101_5 + shifted_state99_105_3 + shifted_state99_105_4 + shifted_state99_105_6 + shifted_state99_105_7 + shifted_state99_106_1 + shifted_state99_106_2 + shifted_state99_109_4 + shifted_state99_116_1 + shifted_state99_118_2 + shifted_state99_118_5 + shifted_state99_118_6 + shifted_state99_118_7 + shifted_state99_132_0 + shifted_state99_132_1 + shifted_state99_132_3 + shifted_state99_132_4 + shifted_state99_132_5 + shifted_state99_132_6 + shifted_state99_132_7 + shifted_state99_133_0 + shifted_state99_133_1 + shifted_state99_133_2 + shifted_state99_133_4 + shifted_state99_133_5 + shifted_state99_133_6 + shifted_state99_133_7 + shifted_state99_141_4 + shifted_state99_141_5 + shifted_state99_141_6 + shifted_state99_141_7 + shifted_state99_142_3 + shifted_state99_142_4 + shifted_state99_142_5 + shifted_state99_142_6 + shifted_state99_142_7 + shifted_state99_152_0 + shifted_state99_152_3 + shifted_state99_156_0 + shifted_state99_156_1 + shifted_state99_156_2 + shifted_state99_156_4 + shifted_state99_181_0 + shifted_state99_181_5 + shifted_state99_181_6 + shifted_state99_181_7 + shifted_state99_187_4 + shifted_state99_197_2 + shifted_state99_197_3 + shifted_state99_197_4 + shifted_state99_197_5);
      reservoir_sum_parallel[100] = (shifted_state100_2_1 + shifted_state100_2_2 + shifted_state100_2_4 + shifted_state100_4_1 + shifted_state100_4_4 + shifted_state100_4_6 + shifted_state100_4_7 + shifted_state100_29_1 + shifted_state100_29_5 + shifted_state100_29_6 + shifted_state100_29_7 + shifted_state100_39_0 + shifted_state100_39_4 + shifted_state100_41_1 + shifted_state100_41_2 + shifted_state100_41_3 + shifted_state100_41_4 + shifted_state100_41_6 + shifted_state100_41_7 + shifted_state100_62_1 + shifted_state100_62_2 + shifted_state100_62_3 + shifted_state100_62_5 + shifted_state100_62_6 + shifted_state100_62_7 + shifted_state100_78_1 + shifted_state100_78_2 + shifted_state100_78_3 + shifted_state100_78_6 + shifted_state100_78_7 + shifted_state100_106_0 + shifted_state100_106_4 + shifted_state100_106_5 + shifted_state100_106_6 + shifted_state100_106_7 + shifted_state100_109_2 + shifted_state100_109_3 + shifted_state100_111_0 + shifted_state100_111_2 + shifted_state100_111_3 + shifted_state100_111_5 + shifted_state100_111_6 + shifted_state100_111_7 + shifted_state100_120_1 + shifted_state100_120_6 + shifted_state100_136_0 + shifted_state100_136_1 + shifted_state100_136_4 + shifted_state100_136_5 + shifted_state100_136_6 + shifted_state100_136_7 + shifted_state100_166_0 + shifted_state100_166_1 + shifted_state100_166_2 + shifted_state100_166_3 + shifted_state100_166_5 + shifted_state100_166_6 + shifted_state100_166_7 + shifted_state100_168_0 + shifted_state100_168_5 + shifted_state100_168_6 + shifted_state100_168_7 + shifted_state100_173_0 + shifted_state100_173_2 + shifted_state100_177_0 + shifted_state100_177_3 + shifted_state100_184_0 + shifted_state100_184_3 + shifted_state100_184_4 + shifted_state100_184_5 + shifted_state100_184_6 + shifted_state100_184_7 + shifted_state100_199_2 + shifted_state100_199_3 + shifted_state100_199_4 + shifted_state100_199_6 + shifted_state100_199_7);
      reservoir_sum_parallel[101] = (shifted_state101_8_0 + shifted_state101_24_4 + shifted_state101_24_5 + shifted_state101_24_6 + shifted_state101_24_7 + shifted_state101_31_0 + shifted_state101_31_1 + shifted_state101_31_3 + shifted_state101_31_4 + shifted_state101_34_0 + shifted_state101_34_3 + shifted_state101_34_4 + shifted_state101_34_5 + shifted_state101_34_6 + shifted_state101_34_7 + shifted_state101_45_0 + shifted_state101_45_1 + shifted_state101_45_3 + shifted_state101_55_1 + shifted_state101_55_5 + shifted_state101_56_1 + shifted_state101_56_3 + shifted_state101_56_5 + shifted_state101_81_0 + shifted_state101_81_1 + shifted_state101_81_2 + shifted_state101_81_3 + shifted_state101_81_4 + shifted_state101_81_5 + shifted_state101_81_6 + shifted_state101_81_7 + shifted_state101_85_1 + shifted_state101_86_0 + shifted_state101_86_1 + shifted_state101_86_2 + shifted_state101_86_4 + shifted_state101_86_5 + shifted_state101_92_0 + shifted_state101_92_1 + shifted_state101_92_5 + shifted_state101_92_6 + shifted_state101_92_7 + shifted_state101_99_3 + shifted_state101_99_4 + shifted_state101_99_5 + shifted_state101_99_6 + shifted_state101_99_7 + shifted_state101_123_1 + shifted_state101_123_2 + shifted_state101_123_4 + shifted_state101_123_5 + shifted_state101_123_6 + shifted_state101_123_7 + shifted_state101_137_0 + shifted_state101_137_1 + shifted_state101_137_3 + shifted_state101_137_5 + shifted_state101_137_6 + shifted_state101_137_7 + shifted_state101_149_3 + shifted_state101_149_4 + shifted_state101_149_6 + shifted_state101_149_7 + shifted_state101_157_1 + shifted_state101_157_4 + shifted_state101_157_6 + shifted_state101_157_7 + shifted_state101_162_3 + shifted_state101_162_4 + shifted_state101_178_0 + shifted_state101_178_4 + shifted_state101_194_0 + shifted_state101_194_4);
      reservoir_sum_parallel[102] = (shifted_state102_5_0 + shifted_state102_5_2 + shifted_state102_16_1 + shifted_state102_16_2 + shifted_state102_16_3 + shifted_state102_16_4 + shifted_state102_16_5 + shifted_state102_16_6 + shifted_state102_16_7 + shifted_state102_17_0 + shifted_state102_17_1 + shifted_state102_17_3 + shifted_state102_17_5 + shifted_state102_17_6 + shifted_state102_17_7 + shifted_state102_25_2 + shifted_state102_25_3 + shifted_state102_25_5 + shifted_state102_25_6 + shifted_state102_25_7 + shifted_state102_31_0 + shifted_state102_31_4 + shifted_state102_36_2 + shifted_state102_36_5 + shifted_state102_36_6 + shifted_state102_36_7 + shifted_state102_37_1 + shifted_state102_37_5 + shifted_state102_40_3 + shifted_state102_45_0 + shifted_state102_45_3 + shifted_state102_45_4 + shifted_state102_45_5 + shifted_state102_45_6 + shifted_state102_45_7 + shifted_state102_57_0 + shifted_state102_57_1 + shifted_state102_57_2 + shifted_state102_57_4 + shifted_state102_89_0 + shifted_state102_89_1 + shifted_state102_89_2 + shifted_state102_89_4 + shifted_state102_89_5 + shifted_state102_89_6 + shifted_state102_89_7 + shifted_state102_102_2 + shifted_state102_102_3 + shifted_state102_102_5 + shifted_state102_102_6 + shifted_state102_102_7 + shifted_state102_111_0 + shifted_state102_111_1 + shifted_state102_111_5 + shifted_state102_111_6 + shifted_state102_111_7 + shifted_state102_120_0 + shifted_state102_120_1 + shifted_state102_120_2 + shifted_state102_130_1 + shifted_state102_130_4 + shifted_state102_133_3 + shifted_state102_133_4 + shifted_state102_135_0 + shifted_state102_135_1 + shifted_state102_135_2 + shifted_state102_135_5 + shifted_state102_135_6 + shifted_state102_135_7 + shifted_state102_146_0 + shifted_state102_146_1 + shifted_state102_146_2 + shifted_state102_146_3 + shifted_state102_146_5 + shifted_state102_146_6 + shifted_state102_146_7 + shifted_state102_164_0 + shifted_state102_164_1 + shifted_state102_164_5 + shifted_state102_164_6 + shifted_state102_164_7 + shifted_state102_171_3 + shifted_state102_171_4 + shifted_state102_171_6 + shifted_state102_174_2 + shifted_state102_198_1 + shifted_state102_198_3);
      reservoir_sum_parallel[103] = (shifted_state103_7_0 + shifted_state103_7_4 + shifted_state103_7_5 + shifted_state103_7_6 + shifted_state103_7_7 + shifted_state103_9_1 + shifted_state103_9_3 + shifted_state103_9_5 + shifted_state103_9_6 + shifted_state103_9_7 + shifted_state103_16_1 + shifted_state103_16_2 + shifted_state103_16_3 + shifted_state103_16_5 + shifted_state103_29_1 + shifted_state103_29_4 + shifted_state103_29_5 + shifted_state103_29_6 + shifted_state103_29_7 + shifted_state103_31_5 + shifted_state103_31_6 + shifted_state103_31_7 + shifted_state103_38_0 + shifted_state103_38_2 + shifted_state103_38_5 + shifted_state103_38_7 + shifted_state103_44_0 + shifted_state103_44_1 + shifted_state103_44_2 + shifted_state103_44_3 + shifted_state103_44_5 + shifted_state103_44_6 + shifted_state103_44_7 + shifted_state103_47_0 + shifted_state103_47_1 + shifted_state103_47_2 + shifted_state103_47_4 + shifted_state103_47_5 + shifted_state103_47_6 + shifted_state103_47_7 + shifted_state103_50_4 + shifted_state103_50_5 + shifted_state103_50_6 + shifted_state103_50_7 + shifted_state103_60_0 + shifted_state103_60_2 + shifted_state103_60_3 + shifted_state103_60_5 + shifted_state103_60_6 + shifted_state103_60_7 + shifted_state103_61_0 + shifted_state103_61_1 + shifted_state103_61_2 + shifted_state103_61_5 + shifted_state103_61_6 + shifted_state103_61_7 + shifted_state103_73_0 + shifted_state103_73_2 + shifted_state103_82_0 + shifted_state103_82_4 + shifted_state103_92_0 + shifted_state103_92_2 + shifted_state103_92_5 + shifted_state103_100_5 + shifted_state103_100_6 + shifted_state103_100_7 + shifted_state103_109_0 + shifted_state103_109_1 + shifted_state103_109_5 + shifted_state103_109_6 + shifted_state103_109_7 + shifted_state103_112_0 + shifted_state103_112_2 + shifted_state103_112_3 + shifted_state103_112_4 + shifted_state103_112_6 + shifted_state103_112_7 + shifted_state103_136_1 + shifted_state103_136_2 + shifted_state103_136_3 + shifted_state103_142_2 + shifted_state103_173_1 + shifted_state103_173_2 + shifted_state103_173_6 + shifted_state103_173_7);
      reservoir_sum_parallel[104] = (shifted_state104_21_0 + shifted_state104_21_1 + shifted_state104_21_3 + shifted_state104_21_4 + shifted_state104_21_6 + shifted_state104_21_7 + shifted_state104_35_1 + shifted_state104_35_3 + shifted_state104_44_0 + shifted_state104_44_3 + shifted_state104_44_5 + shifted_state104_44_6 + shifted_state104_44_7 + shifted_state104_62_0 + shifted_state104_62_1 + shifted_state104_62_5 + shifted_state104_62_6 + shifted_state104_62_7 + shifted_state104_88_0 + shifted_state104_88_1 + shifted_state104_88_3 + shifted_state104_90_0 + shifted_state104_90_2 + shifted_state104_90_4 + shifted_state104_90_5 + shifted_state104_90_6 + shifted_state104_90_7 + shifted_state104_97_1 + shifted_state104_97_4 + shifted_state104_97_6 + shifted_state104_97_7 + shifted_state104_136_0 + shifted_state104_136_2 + shifted_state104_136_4 + shifted_state104_140_0 + shifted_state104_140_2 + shifted_state104_140_4 + shifted_state104_140_5 + shifted_state104_140_6 + shifted_state104_140_7 + shifted_state104_159_2 + shifted_state104_159_3 + shifted_state104_166_0 + shifted_state104_166_1 + shifted_state104_166_3 + shifted_state104_166_4 + shifted_state104_166_5 + shifted_state104_166_7 + shifted_state104_171_1 + shifted_state104_171_2 + shifted_state104_171_5 + shifted_state104_172_0 + shifted_state104_172_1 + shifted_state104_172_3 + shifted_state104_172_5 + shifted_state104_198_5 + shifted_state104_198_6 + shifted_state104_198_7);
      reservoir_sum_parallel[105] = (shifted_state105_1_2 + shifted_state105_1_4 + shifted_state105_1_5 + shifted_state105_1_6 + shifted_state105_1_7 + shifted_state105_2_1 + shifted_state105_2_2 + shifted_state105_2_3 + shifted_state105_2_5 + shifted_state105_2_6 + shifted_state105_2_7 + shifted_state105_25_0 + shifted_state105_25_1 + shifted_state105_25_2 + shifted_state105_25_4 + shifted_state105_25_5 + shifted_state105_25_6 + shifted_state105_25_7 + shifted_state105_30_0 + shifted_state105_30_2 + shifted_state105_42_2 + shifted_state105_42_3 + shifted_state105_53_2 + shifted_state105_53_5 + shifted_state105_57_0 + shifted_state105_57_5 + shifted_state105_57_6 + shifted_state105_57_7 + shifted_state105_59_0 + shifted_state105_59_1 + shifted_state105_59_2 + shifted_state105_59_3 + shifted_state105_59_4 + shifted_state105_59_5 + shifted_state105_59_6 + shifted_state105_59_7 + shifted_state105_62_1 + shifted_state105_62_4 + shifted_state105_62_5 + shifted_state105_62_6 + shifted_state105_62_7 + shifted_state105_70_0 + shifted_state105_70_1 + shifted_state105_70_2 + shifted_state105_70_4 + shifted_state105_70_5 + shifted_state105_70_6 + shifted_state105_70_7 + shifted_state105_87_0 + shifted_state105_87_2 + shifted_state105_87_3 + shifted_state105_87_4 + shifted_state105_87_5 + shifted_state105_87_6 + shifted_state105_87_7 + shifted_state105_91_5 + shifted_state105_99_1 + shifted_state105_99_2 + shifted_state105_99_3 + shifted_state105_99_5 + shifted_state105_99_6 + shifted_state105_99_7 + shifted_state105_102_2 + shifted_state105_102_3 + shifted_state105_102_4 + shifted_state105_105_0 + shifted_state105_105_1 + shifted_state105_105_3 + shifted_state105_105_4 + shifted_state105_105_5 + shifted_state105_110_3 + shifted_state105_110_4 + shifted_state105_110_5 + shifted_state105_110_6 + shifted_state105_110_7 + shifted_state105_112_1 + shifted_state105_112_2 + shifted_state105_112_4 + shifted_state105_118_0 + shifted_state105_118_1 + shifted_state105_118_2 + shifted_state105_118_3 + shifted_state105_118_4 + shifted_state105_118_5 + shifted_state105_118_6 + shifted_state105_118_7 + shifted_state105_120_0 + shifted_state105_120_3 + shifted_state105_120_4 + shifted_state105_130_1 + shifted_state105_130_2 + shifted_state105_130_3 + shifted_state105_130_5 + shifted_state105_139_0 + shifted_state105_139_2 + shifted_state105_139_3 + shifted_state105_139_4 + shifted_state105_139_5 + shifted_state105_139_6 + shifted_state105_139_7 + shifted_state105_149_3 + shifted_state105_149_4 + shifted_state105_154_1 + shifted_state105_154_2 + shifted_state105_154_4 + shifted_state105_154_6 + shifted_state105_154_7 + shifted_state105_160_3 + shifted_state105_190_0 + shifted_state105_190_1 + shifted_state105_190_4);
      reservoir_sum_parallel[106] = (shifted_state106_10_0 + shifted_state106_10_1 + shifted_state106_10_5 + shifted_state106_10_6 + shifted_state106_10_7 + shifted_state106_21_0 + shifted_state106_21_1 + shifted_state106_21_2 + shifted_state106_21_3 + shifted_state106_21_5 + shifted_state106_21_6 + shifted_state106_21_7 + shifted_state106_23_4 + shifted_state106_23_6 + shifted_state106_23_7 + shifted_state106_35_1 + shifted_state106_35_2 + shifted_state106_35_4 + shifted_state106_35_5 + shifted_state106_52_1 + shifted_state106_52_2 + shifted_state106_52_3 + shifted_state106_52_5 + shifted_state106_52_6 + shifted_state106_52_7 + shifted_state106_59_1 + shifted_state106_59_2 + shifted_state106_59_5 + shifted_state106_59_6 + shifted_state106_59_7 + shifted_state106_62_1 + shifted_state106_62_3 + shifted_state106_85_1 + shifted_state106_85_2 + shifted_state106_85_4 + shifted_state106_85_5 + shifted_state106_96_1 + shifted_state106_96_2 + shifted_state106_96_3 + shifted_state106_96_6 + shifted_state106_96_7 + shifted_state106_114_0 + shifted_state106_114_5 + shifted_state106_114_6 + shifted_state106_114_7 + shifted_state106_120_1 + shifted_state106_120_4 + shifted_state106_126_5 + shifted_state106_138_2 + shifted_state106_138_5 + shifted_state106_138_6 + shifted_state106_138_7 + shifted_state106_144_0 + shifted_state106_144_2 + shifted_state106_144_3 + shifted_state106_144_4 + shifted_state106_151_0 + shifted_state106_151_3 + shifted_state106_151_6 + shifted_state106_151_7 + shifted_state106_179_0 + shifted_state106_179_1 + shifted_state106_179_4 + shifted_state106_179_5 + shifted_state106_179_6 + shifted_state106_179_7 + shifted_state106_198_0 + shifted_state106_198_6 + shifted_state106_199_2 + shifted_state106_199_3 + shifted_state106_199_4);
      reservoir_sum_parallel[107] = (shifted_state107_5_1 + shifted_state107_5_2 + shifted_state107_5_4 + shifted_state107_6_0 + shifted_state107_6_2 + shifted_state107_21_1 + shifted_state107_21_4 + shifted_state107_21_5 + shifted_state107_21_6 + shifted_state107_21_7 + shifted_state107_35_0 + shifted_state107_35_3 + shifted_state107_35_4 + shifted_state107_48_0 + shifted_state107_48_1 + shifted_state107_48_2 + shifted_state107_48_3 + shifted_state107_48_4 + shifted_state107_48_5 + shifted_state107_48_7 + shifted_state107_49_2 + shifted_state107_49_3 + shifted_state107_75_0 + shifted_state107_75_3 + shifted_state107_82_0 + shifted_state107_82_3 + shifted_state107_82_4 + shifted_state107_88_0 + shifted_state107_88_1 + shifted_state107_120_0 + shifted_state107_120_2 + shifted_state107_120_3 + shifted_state107_120_4 + shifted_state107_120_5 + shifted_state107_120_6 + shifted_state107_120_7 + shifted_state107_133_0 + shifted_state107_133_3 + shifted_state107_148_0 + shifted_state107_148_1 + shifted_state107_148_3 + shifted_state107_184_1 + shifted_state107_184_3 + shifted_state107_184_4 + shifted_state107_184_5 + shifted_state107_184_6 + shifted_state107_184_7);
      reservoir_sum_parallel[108] = (shifted_state108_14_5 + shifted_state108_15_0 + shifted_state108_15_1 + shifted_state108_15_3 + shifted_state108_18_0 + shifted_state108_18_4 + shifted_state108_19_0 + shifted_state108_19_1 + shifted_state108_19_4 + shifted_state108_19_5 + shifted_state108_19_6 + shifted_state108_19_7 + shifted_state108_32_2 + shifted_state108_32_3 + shifted_state108_32_4 + shifted_state108_36_0 + shifted_state108_36_2 + shifted_state108_39_0 + shifted_state108_39_1 + shifted_state108_39_3 + shifted_state108_41_0 + shifted_state108_41_1 + shifted_state108_41_4 + shifted_state108_62_0 + shifted_state108_62_2 + shifted_state108_62_5 + shifted_state108_62_6 + shifted_state108_62_7 + shifted_state108_67_2 + shifted_state108_67_5 + shifted_state108_67_6 + shifted_state108_67_7 + shifted_state108_77_0 + shifted_state108_77_1 + shifted_state108_81_0 + shifted_state108_81_3 + shifted_state108_91_1 + shifted_state108_91_4 + shifted_state108_91_5 + shifted_state108_91_6 + shifted_state108_91_7 + shifted_state108_97_0 + shifted_state108_97_1 + shifted_state108_97_2 + shifted_state108_97_4 + shifted_state108_97_5 + shifted_state108_97_6 + shifted_state108_97_7 + shifted_state108_98_0 + shifted_state108_98_4 + shifted_state108_130_1 + shifted_state108_130_4 + shifted_state108_130_5 + shifted_state108_130_6 + shifted_state108_130_7 + shifted_state108_132_2 + shifted_state108_132_3 + shifted_state108_132_4 + shifted_state108_132_5 + shifted_state108_132_6 + shifted_state108_132_7 + shifted_state108_151_1 + shifted_state108_151_2 + shifted_state108_151_3 + shifted_state108_151_6 + shifted_state108_151_7 + shifted_state108_159_1 + shifted_state108_159_3 + shifted_state108_159_5 + shifted_state108_159_6 + shifted_state108_159_7 + shifted_state108_173_1 + shifted_state108_173_2 + shifted_state108_173_3 + shifted_state108_173_4 + shifted_state108_173_5 + shifted_state108_173_6 + shifted_state108_173_7 + shifted_state108_182_0 + shifted_state108_182_1 + shifted_state108_182_2 + shifted_state108_198_0 + shifted_state108_198_2 + shifted_state108_198_5 + shifted_state108_198_6 + shifted_state108_198_7);
      reservoir_sum_parallel[109] = (shifted_state109_1_0 + shifted_state109_1_2 + shifted_state109_1_3 + shifted_state109_1_4 + shifted_state109_1_5 + shifted_state109_1_6 + shifted_state109_1_7 + shifted_state109_13_0 + shifted_state109_13_3 + shifted_state109_13_4 + shifted_state109_13_5 + shifted_state109_19_3 + shifted_state109_19_4 + shifted_state109_19_5 + shifted_state109_19_6 + shifted_state109_19_7 + shifted_state109_32_0 + shifted_state109_32_2 + shifted_state109_32_3 + shifted_state109_51_3 + shifted_state109_55_1 + shifted_state109_55_2 + shifted_state109_55_3 + shifted_state109_83_0 + shifted_state109_83_4 + shifted_state109_90_2 + shifted_state109_90_3 + shifted_state109_90_4 + shifted_state109_90_5 + shifted_state109_90_6 + shifted_state109_90_7 + shifted_state109_100_0 + shifted_state109_100_4 + shifted_state109_100_5 + shifted_state109_152_2 + shifted_state109_152_3 + shifted_state109_152_5 + shifted_state109_152_6 + shifted_state109_152_7 + shifted_state109_155_1 + shifted_state109_155_3 + shifted_state109_155_5 + shifted_state109_155_6 + shifted_state109_155_7 + shifted_state109_160_3 + shifted_state109_160_5 + shifted_state109_170_0 + shifted_state109_170_1 + shifted_state109_170_2 + shifted_state109_173_1 + shifted_state109_173_2 + shifted_state109_173_4 + shifted_state109_173_6 + shifted_state109_173_7 + shifted_state109_174_0 + shifted_state109_174_2 + shifted_state109_174_5 + shifted_state109_174_6 + shifted_state109_174_7 + shifted_state109_187_0 + shifted_state109_187_1 + shifted_state109_187_5 + shifted_state109_187_6 + shifted_state109_187_7 + shifted_state109_188_2 + shifted_state109_188_5 + shifted_state109_188_6 + shifted_state109_188_7 + shifted_state109_191_0 + shifted_state109_191_1 + shifted_state109_191_2 + shifted_state109_191_5 + shifted_state109_191_6 + shifted_state109_191_7);
      reservoir_sum_parallel[110] = (shifted_state110_11_2 + shifted_state110_11_5 + shifted_state110_15_0 + shifted_state110_15_2 + shifted_state110_15_3 + shifted_state110_15_4 + shifted_state110_30_0 + shifted_state110_30_1 + shifted_state110_30_5 + shifted_state110_53_0 + shifted_state110_53_2 + shifted_state110_53_4 + shifted_state110_53_6 + shifted_state110_53_7 + shifted_state110_58_1 + shifted_state110_58_4 + shifted_state110_59_0 + shifted_state110_59_1 + shifted_state110_59_3 + shifted_state110_59_4 + shifted_state110_59_5 + shifted_state110_59_6 + shifted_state110_59_7 + shifted_state110_65_1 + shifted_state110_65_4 + shifted_state110_68_1 + shifted_state110_68_2 + shifted_state110_68_5 + shifted_state110_70_1 + shifted_state110_70_3 + shifted_state110_70_4 + shifted_state110_70_5 + shifted_state110_70_6 + shifted_state110_70_7 + shifted_state110_76_1 + shifted_state110_76_2 + shifted_state110_76_3 + shifted_state110_76_5 + shifted_state110_76_6 + shifted_state110_76_7 + shifted_state110_85_3 + shifted_state110_85_4 + shifted_state110_114_2 + shifted_state110_114_3 + shifted_state110_114_6 + shifted_state110_114_7 + shifted_state110_124_0 + shifted_state110_124_1 + shifted_state110_124_4 + shifted_state110_129_2 + shifted_state110_129_3 + shifted_state110_129_5 + shifted_state110_138_1 + shifted_state110_138_3 + shifted_state110_138_4 + shifted_state110_138_5 + shifted_state110_138_6 + shifted_state110_138_7 + shifted_state110_147_0 + shifted_state110_147_2 + shifted_state110_147_4 + shifted_state110_155_1 + shifted_state110_155_5 + shifted_state110_158_1 + shifted_state110_158_2 + shifted_state110_161_0 + shifted_state110_161_2 + shifted_state110_161_4 + shifted_state110_165_1 + shifted_state110_165_4 + shifted_state110_165_5 + shifted_state110_171_1 + shifted_state110_171_2 + shifted_state110_171_3 + shifted_state110_171_6 + shifted_state110_171_7 + shifted_state110_172_0 + shifted_state110_172_4 + shifted_state110_174_2 + shifted_state110_174_6 + shifted_state110_174_7 + shifted_state110_179_2 + shifted_state110_179_4 + shifted_state110_179_5 + shifted_state110_179_6 + shifted_state110_179_7 + shifted_state110_181_2 + shifted_state110_181_4 + shifted_state110_181_5 + shifted_state110_181_6 + shifted_state110_181_7 + shifted_state110_193_1 + shifted_state110_193_2 + shifted_state110_199_1 + shifted_state110_199_2 + shifted_state110_199_5 + shifted_state110_199_6 + shifted_state110_199_7);
      reservoir_sum_parallel[111] = (shifted_state111_15_1 + shifted_state111_15_2 + shifted_state111_17_0 + shifted_state111_17_1 + shifted_state111_17_2 + shifted_state111_17_5 + shifted_state111_17_6 + shifted_state111_17_7 + shifted_state111_22_1 + shifted_state111_22_3 + shifted_state111_22_4 + shifted_state111_22_5 + shifted_state111_28_0 + shifted_state111_84_3 + shifted_state111_84_4 + shifted_state111_90_3 + shifted_state111_90_4 + shifted_state111_90_5 + shifted_state111_90_6 + shifted_state111_90_7 + shifted_state111_93_0 + shifted_state111_93_3 + shifted_state111_93_4 + shifted_state111_93_6 + shifted_state111_93_7 + shifted_state111_113_0 + shifted_state111_113_5 + shifted_state111_122_0 + shifted_state111_122_3 + shifted_state111_122_4 + shifted_state111_122_5 + shifted_state111_122_6 + shifted_state111_122_7 + shifted_state111_130_0 + shifted_state111_130_1 + shifted_state111_134_1 + shifted_state111_134_2 + shifted_state111_134_4 + shifted_state111_139_4 + shifted_state111_165_0 + shifted_state111_165_2 + shifted_state111_165_3 + shifted_state111_165_4 + shifted_state111_165_6 + shifted_state111_165_7 + shifted_state111_169_1 + shifted_state111_169_2 + shifted_state111_169_3 + shifted_state111_169_4 + shifted_state111_169_5 + shifted_state111_169_6 + shifted_state111_169_7 + shifted_state111_170_1 + shifted_state111_170_2 + shifted_state111_170_3 + shifted_state111_170_4 + shifted_state111_170_6 + shifted_state111_170_7);
      reservoir_sum_parallel[112] = (shifted_state112_28_2 + shifted_state112_28_3 + shifted_state112_34_1 + shifted_state112_34_2 + shifted_state112_34_3 + shifted_state112_43_3 + shifted_state112_43_4 + shifted_state112_63_0 + shifted_state112_63_1 + shifted_state112_63_2 + shifted_state112_63_3 + shifted_state112_65_0 + shifted_state112_65_1 + shifted_state112_65_5 + shifted_state112_65_6 + shifted_state112_65_7 + shifted_state112_68_0 + shifted_state112_68_1 + shifted_state112_68_3 + shifted_state112_68_4 + shifted_state112_68_5 + shifted_state112_68_6 + shifted_state112_68_7 + shifted_state112_92_0 + shifted_state112_92_1 + shifted_state112_92_2 + shifted_state112_92_3 + shifted_state112_92_4 + shifted_state112_119_1 + shifted_state112_119_4 + shifted_state112_123_4 + shifted_state112_123_5 + shifted_state112_123_6 + shifted_state112_123_7 + shifted_state112_124_0 + shifted_state112_124_5 + shifted_state112_133_0 + shifted_state112_133_1 + shifted_state112_133_3 + shifted_state112_135_0 + shifted_state112_135_4 + shifted_state112_135_5 + shifted_state112_135_6 + shifted_state112_135_7 + shifted_state112_138_4 + shifted_state112_138_5 + shifted_state112_138_6 + shifted_state112_138_7 + shifted_state112_141_0 + shifted_state112_141_3 + shifted_state112_141_6 + shifted_state112_141_7 + shifted_state112_173_0 + shifted_state112_173_1 + shifted_state112_173_2 + shifted_state112_173_3 + shifted_state112_173_4 + shifted_state112_183_0 + shifted_state112_183_1 + shifted_state112_183_4 + shifted_state112_183_5 + shifted_state112_183_7);
      reservoir_sum_parallel[113] = (shifted_state113_10_1 + shifted_state113_10_3 + shifted_state113_24_0 + shifted_state113_24_2 + shifted_state113_24_3 + shifted_state113_24_4 + shifted_state113_31_0 + shifted_state113_31_3 + shifted_state113_31_4 + shifted_state113_31_6 + shifted_state113_31_7 + shifted_state113_32_1 + shifted_state113_32_2 + shifted_state113_32_3 + shifted_state113_36_6 + shifted_state113_36_7 + shifted_state113_40_0 + shifted_state113_40_5 + shifted_state113_54_0 + shifted_state113_54_1 + shifted_state113_54_2 + shifted_state113_54_3 + shifted_state113_54_5 + shifted_state113_77_0 + shifted_state113_77_1 + shifted_state113_77_2 + shifted_state113_84_1 + shifted_state113_84_2 + shifted_state113_84_4 + shifted_state113_84_6 + shifted_state113_84_7 + shifted_state113_87_3 + shifted_state113_87_4 + shifted_state113_95_1 + shifted_state113_95_2 + shifted_state113_95_3 + shifted_state113_95_6 + shifted_state113_95_7 + shifted_state113_105_0 + shifted_state113_105_1 + shifted_state113_105_3 + shifted_state113_105_4 + shifted_state113_105_5 + shifted_state113_105_6 + shifted_state113_105_7 + shifted_state113_123_2 + shifted_state113_123_4 + shifted_state113_123_5 + shifted_state113_136_0 + shifted_state113_136_2 + shifted_state113_136_3 + shifted_state113_136_5 + shifted_state113_136_6 + shifted_state113_136_7 + shifted_state113_148_0 + shifted_state113_148_3 + shifted_state113_152_1 + shifted_state113_152_3 + shifted_state113_152_4 + shifted_state113_152_5 + shifted_state113_152_6 + shifted_state113_152_7 + shifted_state113_174_1 + shifted_state113_174_2 + shifted_state113_174_4 + shifted_state113_188_0 + shifted_state113_188_1 + shifted_state113_188_3 + shifted_state113_188_4 + shifted_state113_198_1 + shifted_state113_198_2 + shifted_state113_198_3 + shifted_state113_198_4 + shifted_state113_198_5 + shifted_state113_198_7);
      reservoir_sum_parallel[114] = (shifted_state114_2_1 + shifted_state114_2_5 + shifted_state114_2_6 + shifted_state114_2_7 + shifted_state114_5_0 + shifted_state114_5_1 + shifted_state114_5_3 + shifted_state114_5_4 + shifted_state114_5_6 + shifted_state114_5_7 + shifted_state114_6_2 + shifted_state114_6_4 + shifted_state114_6_5 + shifted_state114_6_6 + shifted_state114_6_7 + shifted_state114_23_1 + shifted_state114_23_2 + shifted_state114_29_0 + shifted_state114_29_1 + shifted_state114_29_4 + shifted_state114_29_5 + shifted_state114_29_6 + shifted_state114_29_7 + shifted_state114_35_1 + shifted_state114_35_5 + shifted_state114_35_6 + shifted_state114_35_7 + shifted_state114_39_0 + shifted_state114_39_1 + shifted_state114_39_4 + shifted_state114_39_5 + shifted_state114_39_6 + shifted_state114_39_7 + shifted_state114_43_5 + shifted_state114_54_0 + shifted_state114_54_1 + shifted_state114_54_2 + shifted_state114_54_5 + shifted_state114_54_6 + shifted_state114_54_7 + shifted_state114_58_1 + shifted_state114_58_2 + shifted_state114_58_3 + shifted_state114_58_6 + shifted_state114_58_7 + shifted_state114_97_0 + shifted_state114_97_1 + shifted_state114_97_2 + shifted_state114_97_4 + shifted_state114_97_6 + shifted_state114_97_7 + shifted_state114_108_0 + shifted_state114_108_1 + shifted_state114_108_3 + shifted_state114_108_4 + shifted_state114_108_5 + shifted_state114_108_6 + shifted_state114_108_7 + shifted_state114_110_2 + shifted_state114_110_3 + shifted_state114_110_4 + shifted_state114_118_0 + shifted_state114_118_2 + shifted_state114_118_5 + shifted_state114_118_6 + shifted_state114_118_7 + shifted_state114_126_2 + shifted_state114_126_3 + shifted_state114_164_3 + shifted_state114_164_4 + shifted_state114_198_1 + shifted_state114_198_4 + shifted_state114_199_1 + shifted_state114_199_3 + shifted_state114_199_5 + shifted_state114_199_6 + shifted_state114_199_7);
      reservoir_sum_parallel[115] = (shifted_state115_5_1 + shifted_state115_5_2 + shifted_state115_10_0 + shifted_state115_10_1 + shifted_state115_10_4 + shifted_state115_10_5 + shifted_state115_10_6 + shifted_state115_10_7 + shifted_state115_16_0 + shifted_state115_16_1 + shifted_state115_16_4 + shifted_state115_22_1 + shifted_state115_22_2 + shifted_state115_22_5 + shifted_state115_26_3 + shifted_state115_26_5 + shifted_state115_26_6 + shifted_state115_26_7 + shifted_state115_37_4 + shifted_state115_37_5 + shifted_state115_37_6 + shifted_state115_37_7 + shifted_state115_43_0 + shifted_state115_43_4 + shifted_state115_62_1 + shifted_state115_62_2 + shifted_state115_62_4 + shifted_state115_62_6 + shifted_state115_62_7 + shifted_state115_68_0 + shifted_state115_68_6 + shifted_state115_71_0 + shifted_state115_71_2 + shifted_state115_71_5 + shifted_state115_71_6 + shifted_state115_71_7 + shifted_state115_80_6 + shifted_state115_80_7 + shifted_state115_83_1 + shifted_state115_83_3 + shifted_state115_83_4 + shifted_state115_83_5 + shifted_state115_83_6 + shifted_state115_83_7 + shifted_state115_88_1 + shifted_state115_88_2 + shifted_state115_88_5 + shifted_state115_88_6 + shifted_state115_88_7 + shifted_state115_101_0 + shifted_state115_101_1 + shifted_state115_101_2 + shifted_state115_101_4 + shifted_state115_101_5 + shifted_state115_101_6 + shifted_state115_101_7 + shifted_state115_107_0 + shifted_state115_107_1 + shifted_state115_107_2 + shifted_state115_107_3 + shifted_state115_107_4 + shifted_state115_107_5 + shifted_state115_138_0 + shifted_state115_138_6 + shifted_state115_163_0 + shifted_state115_163_1 + shifted_state115_163_3 + shifted_state115_171_2 + shifted_state115_171_3 + shifted_state115_171_4 + shifted_state115_175_0 + shifted_state115_175_2 + shifted_state115_175_5 + shifted_state115_175_6 + shifted_state115_175_7 + shifted_state115_176_0 + shifted_state115_176_1 + shifted_state115_176_2 + shifted_state115_176_4 + shifted_state115_176_5 + shifted_state115_176_6 + shifted_state115_176_7 + shifted_state115_178_1 + shifted_state115_178_3 + shifted_state115_178_4 + shifted_state115_179_0 + shifted_state115_179_1 + shifted_state115_179_5 + shifted_state115_185_0 + shifted_state115_185_1 + shifted_state115_185_4 + shifted_state115_191_2 + shifted_state115_191_3 + shifted_state115_191_4 + shifted_state115_191_6 + shifted_state115_191_7 + shifted_state115_199_1 + shifted_state115_199_2 + shifted_state115_199_3 + shifted_state115_199_5);
      reservoir_sum_parallel[116] = (shifted_state116_3_0 + shifted_state116_3_2 + shifted_state116_3_3 + shifted_state116_3_4 + shifted_state116_3_6 + shifted_state116_3_7 + shifted_state116_10_0 + shifted_state116_10_1 + shifted_state116_10_3 + shifted_state116_10_4 + shifted_state116_10_6 + shifted_state116_10_7 + shifted_state116_23_0 + shifted_state116_23_1 + shifted_state116_23_3 + shifted_state116_23_6 + shifted_state116_26_1 + shifted_state116_26_4 + shifted_state116_26_5 + shifted_state116_26_6 + shifted_state116_26_7 + shifted_state116_28_0 + shifted_state116_28_1 + shifted_state116_28_2 + shifted_state116_28_3 + shifted_state116_28_4 + shifted_state116_29_0 + shifted_state116_29_2 + shifted_state116_29_3 + shifted_state116_29_4 + shifted_state116_71_0 + shifted_state116_71_3 + shifted_state116_71_4 + shifted_state116_72_4 + shifted_state116_72_6 + shifted_state116_72_7 + shifted_state116_73_3 + shifted_state116_73_4 + shifted_state116_80_4 + shifted_state116_80_6 + shifted_state116_80_7 + shifted_state116_83_0 + shifted_state116_83_1 + shifted_state116_83_2 + shifted_state116_83_3 + shifted_state116_83_4 + shifted_state116_83_5 + shifted_state116_83_6 + shifted_state116_83_7 + shifted_state116_91_4 + shifted_state116_112_1 + shifted_state116_112_2 + shifted_state116_112_4 + shifted_state116_112_6 + shifted_state116_112_7 + shifted_state116_122_0 + shifted_state116_139_1 + shifted_state116_139_2 + shifted_state116_139_6 + shifted_state116_139_7 + shifted_state116_140_1 + shifted_state116_140_2 + shifted_state116_140_5 + shifted_state116_152_0 + shifted_state116_152_3 + shifted_state116_152_4 + shifted_state116_152_5 + shifted_state116_153_6 + shifted_state116_154_0 + shifted_state116_154_1 + shifted_state116_154_3 + shifted_state116_154_4 + shifted_state116_154_5 + shifted_state116_155_0 + shifted_state116_155_1 + shifted_state116_155_2 + shifted_state116_155_3 + shifted_state116_155_4 + shifted_state116_155_5 + shifted_state116_155_6 + shifted_state116_155_7 + shifted_state116_161_1 + shifted_state116_161_4 + shifted_state116_161_5 + shifted_state116_161_6 + shifted_state116_161_7 + shifted_state116_175_3 + shifted_state116_175_5 + shifted_state116_175_6 + shifted_state116_175_7);
      reservoir_sum_parallel[117] = (shifted_state117_4_2 + shifted_state117_4_5 + shifted_state117_4_6 + shifted_state117_4_7 + shifted_state117_7_0 + shifted_state117_7_1 + shifted_state117_7_2 + shifted_state117_16_0 + shifted_state117_16_2 + shifted_state117_16_5 + shifted_state117_36_0 + shifted_state117_36_2 + shifted_state117_36_3 + shifted_state117_36_4 + shifted_state117_45_0 + shifted_state117_45_1 + shifted_state117_45_5 + shifted_state117_45_6 + shifted_state117_45_7 + shifted_state117_68_2 + shifted_state117_68_3 + shifted_state117_68_5 + shifted_state117_68_6 + shifted_state117_68_7 + shifted_state117_72_2 + shifted_state117_72_5 + shifted_state117_77_0 + shifted_state117_77_2 + shifted_state117_77_3 + shifted_state117_77_6 + shifted_state117_77_7 + shifted_state117_81_1 + shifted_state117_81_4 + shifted_state117_81_5 + shifted_state117_81_6 + shifted_state117_81_7 + shifted_state117_101_1 + shifted_state117_101_2 + shifted_state117_101_3 + shifted_state117_124_0 + shifted_state117_132_0 + shifted_state117_141_2 + shifted_state117_141_4 + shifted_state117_141_5 + shifted_state117_141_6 + shifted_state117_141_7 + shifted_state117_144_1 + shifted_state117_144_3 + shifted_state117_144_4 + shifted_state117_144_5 + shifted_state117_144_6 + shifted_state117_144_7 + shifted_state117_152_0 + shifted_state117_152_3 + shifted_state117_152_4 + shifted_state117_152_5 + shifted_state117_152_6 + shifted_state117_152_7 + shifted_state117_163_0 + shifted_state117_163_1 + shifted_state117_163_3 + shifted_state117_163_5 + shifted_state117_163_6 + shifted_state117_163_7 + shifted_state117_193_3 + shifted_state117_193_6 + shifted_state117_193_7);
      reservoir_sum_parallel[118] = (shifted_state118_1_0 + shifted_state118_1_3 + shifted_state118_1_4 + shifted_state118_1_5 + shifted_state118_1_6 + shifted_state118_1_7 + shifted_state118_6_1 + shifted_state118_6_4 + shifted_state118_6_5 + shifted_state118_6_6 + shifted_state118_6_7 + shifted_state118_9_0 + shifted_state118_9_1 + shifted_state118_9_3 + shifted_state118_9_5 + shifted_state118_9_6 + shifted_state118_9_7 + shifted_state118_11_0 + shifted_state118_11_1 + shifted_state118_11_4 + shifted_state118_11_5 + shifted_state118_11_6 + shifted_state118_11_7 + shifted_state118_20_1 + shifted_state118_20_3 + shifted_state118_20_4 + shifted_state118_20_5 + shifted_state118_20_6 + shifted_state118_20_7 + shifted_state118_25_0 + shifted_state118_25_2 + shifted_state118_25_4 + shifted_state118_28_2 + shifted_state118_28_5 + shifted_state118_28_6 + shifted_state118_28_7 + shifted_state118_65_0 + shifted_state118_65_1 + shifted_state118_65_2 + shifted_state118_74_1 + shifted_state118_74_4 + shifted_state118_74_5 + shifted_state118_79_3 + shifted_state118_85_1 + shifted_state118_85_2 + shifted_state118_85_5 + shifted_state118_85_6 + shifted_state118_85_7 + shifted_state118_88_0 + shifted_state118_88_1 + shifted_state118_88_2 + shifted_state118_100_0 + shifted_state118_100_4 + shifted_state118_100_5 + shifted_state118_100_6 + shifted_state118_100_7 + shifted_state118_115_0 + shifted_state118_115_1 + shifted_state118_115_2 + shifted_state118_122_3 + shifted_state118_122_5 + shifted_state118_122_6 + shifted_state118_122_7 + shifted_state118_139_0 + shifted_state118_139_3 + shifted_state118_139_6 + shifted_state118_147_2 + shifted_state118_147_5 + shifted_state118_147_6 + shifted_state118_147_7 + shifted_state118_158_1 + shifted_state118_190_0 + shifted_state118_190_1 + shifted_state118_190_3);
      reservoir_sum_parallel[119] = (shifted_state119_3_1 + shifted_state119_3_4 + shifted_state119_3_5 + shifted_state119_3_6 + shifted_state119_3_7 + shifted_state119_7_4 + shifted_state119_7_5 + shifted_state119_7_7 + shifted_state119_26_0 + shifted_state119_26_1 + shifted_state119_26_3 + shifted_state119_26_4 + shifted_state119_26_5 + shifted_state119_26_6 + shifted_state119_26_7 + shifted_state119_51_0 + shifted_state119_51_1 + shifted_state119_51_2 + shifted_state119_51_5 + shifted_state119_51_6 + shifted_state119_51_7 + shifted_state119_53_4 + shifted_state119_53_5 + shifted_state119_53_6 + shifted_state119_53_7 + shifted_state119_56_1 + shifted_state119_56_2 + shifted_state119_56_5 + shifted_state119_56_6 + shifted_state119_56_7 + shifted_state119_57_1 + shifted_state119_57_4 + shifted_state119_57_5 + shifted_state119_57_6 + shifted_state119_57_7 + shifted_state119_69_0 + shifted_state119_95_0 + shifted_state119_95_2 + shifted_state119_95_3 + shifted_state119_95_4 + shifted_state119_95_5 + shifted_state119_95_6 + shifted_state119_95_7 + shifted_state119_103_4 + shifted_state119_114_0 + shifted_state119_124_0 + shifted_state119_124_5 + shifted_state119_124_6 + shifted_state119_124_7 + shifted_state119_130_0 + shifted_state119_130_1 + shifted_state119_130_2 + shifted_state119_130_4 + shifted_state119_144_1 + shifted_state119_144_2 + shifted_state119_144_3 + shifted_state119_167_3 + shifted_state119_167_5 + shifted_state119_167_6 + shifted_state119_167_7 + shifted_state119_168_0 + shifted_state119_168_2 + shifted_state119_168_3 + shifted_state119_168_4 + shifted_state119_192_0 + shifted_state119_192_1 + shifted_state119_192_2 + shifted_state119_192_3 + shifted_state119_192_4 + shifted_state119_192_5 + shifted_state119_192_6 + shifted_state119_192_7);
      reservoir_sum_parallel[120] = (shifted_state120_2_2 + shifted_state120_2_3 + shifted_state120_2_5 + shifted_state120_2_6 + shifted_state120_2_7 + shifted_state120_21_0 + shifted_state120_21_1 + shifted_state120_21_2 + shifted_state120_21_3 + shifted_state120_21_4 + shifted_state120_21_5 + shifted_state120_21_6 + shifted_state120_21_7 + shifted_state120_31_0 + shifted_state120_31_2 + shifted_state120_31_3 + shifted_state120_37_0 + shifted_state120_37_1 + shifted_state120_48_4 + shifted_state120_57_1 + shifted_state120_57_2 + shifted_state120_57_4 + shifted_state120_57_5 + shifted_state120_57_6 + shifted_state120_57_7 + shifted_state120_70_1 + shifted_state120_70_2 + shifted_state120_70_3 + shifted_state120_70_5 + shifted_state120_70_6 + shifted_state120_70_7 + shifted_state120_74_1 + shifted_state120_74_3 + shifted_state120_74_4 + shifted_state120_76_1 + shifted_state120_76_3 + shifted_state120_76_5 + shifted_state120_98_0 + shifted_state120_98_1 + shifted_state120_98_2 + shifted_state120_98_3 + shifted_state120_98_4 + shifted_state120_98_5 + shifted_state120_98_6 + shifted_state120_98_7 + shifted_state120_124_0 + shifted_state120_124_1 + shifted_state120_124_2 + shifted_state120_124_4 + shifted_state120_124_5 + shifted_state120_124_6 + shifted_state120_124_7 + shifted_state120_162_1 + shifted_state120_162_3 + shifted_state120_162_4 + shifted_state120_164_0 + shifted_state120_164_1 + shifted_state120_171_0 + shifted_state120_171_1 + shifted_state120_171_2 + shifted_state120_171_3 + shifted_state120_171_5 + shifted_state120_171_6 + shifted_state120_171_7 + shifted_state120_180_0 + shifted_state120_180_1 + shifted_state120_180_3 + shifted_state120_180_4 + shifted_state120_180_5 + shifted_state120_180_6 + shifted_state120_180_7 + shifted_state120_182_0 + shifted_state120_182_2 + shifted_state120_182_3 + shifted_state120_182_4);
      reservoir_sum_parallel[121] = (shifted_state121_14_0 + shifted_state121_14_1 + shifted_state121_14_3 + shifted_state121_14_5 + shifted_state121_28_1 + shifted_state121_28_4 + shifted_state121_28_6 + shifted_state121_28_7 + shifted_state121_70_0 + shifted_state121_70_2 + shifted_state121_70_3 + shifted_state121_72_1 + shifted_state121_72_5 + shifted_state121_82_0 + shifted_state121_82_1 + shifted_state121_82_2 + shifted_state121_82_4 + shifted_state121_82_5 + shifted_state121_82_6 + shifted_state121_82_7 + shifted_state121_86_0 + shifted_state121_86_1 + shifted_state121_86_2 + shifted_state121_86_5 + shifted_state121_101_1 + shifted_state121_101_4 + shifted_state121_101_5 + shifted_state121_101_6 + shifted_state121_101_7 + shifted_state121_133_0 + shifted_state121_133_2 + shifted_state121_133_3 + shifted_state121_133_5 + shifted_state121_185_0 + shifted_state121_185_3 + shifted_state121_185_4 + shifted_state121_185_6 + shifted_state121_185_7 + shifted_state121_187_0 + shifted_state121_187_1 + shifted_state121_187_2 + shifted_state121_187_3 + shifted_state121_187_5 + shifted_state121_187_7);
      reservoir_sum_parallel[122] = (shifted_state122_16_0 + shifted_state122_16_2 + shifted_state122_16_4 + shifted_state122_16_5 + shifted_state122_16_6 + shifted_state122_16_7 + shifted_state122_17_1 + shifted_state122_17_2 + shifted_state122_17_5 + shifted_state122_17_6 + shifted_state122_17_7 + shifted_state122_18_0 + shifted_state122_18_2 + shifted_state122_18_5 + shifted_state122_18_6 + shifted_state122_18_7 + shifted_state122_21_0 + shifted_state122_21_1 + shifted_state122_21_4 + shifted_state122_21_6 + shifted_state122_21_7 + shifted_state122_22_0 + shifted_state122_22_1 + shifted_state122_22_2 + shifted_state122_22_3 + shifted_state122_22_6 + shifted_state122_23_1 + shifted_state122_45_1 + shifted_state122_45_3 + shifted_state122_45_4 + shifted_state122_45_6 + shifted_state122_45_7 + shifted_state122_55_2 + shifted_state122_55_4 + shifted_state122_55_6 + shifted_state122_55_7 + shifted_state122_90_2 + shifted_state122_90_3 + shifted_state122_91_2 + shifted_state122_91_3 + shifted_state122_91_5 + shifted_state122_91_6 + shifted_state122_91_7 + shifted_state122_94_0 + shifted_state122_94_3 + shifted_state122_97_5 + shifted_state122_97_6 + shifted_state122_97_7 + shifted_state122_112_1 + shifted_state122_112_2 + shifted_state122_112_3 + shifted_state122_114_2 + shifted_state122_114_4 + shifted_state122_114_6 + shifted_state122_114_7 + shifted_state122_142_2 + shifted_state122_142_5 + shifted_state122_143_0 + shifted_state122_143_3 + shifted_state122_143_4 + shifted_state122_143_5 + shifted_state122_143_6 + shifted_state122_143_7 + shifted_state122_154_2 + shifted_state122_154_5 + shifted_state122_154_6 + shifted_state122_154_7 + shifted_state122_175_0 + shifted_state122_175_1 + shifted_state122_175_5 + shifted_state122_182_0 + shifted_state122_182_1 + shifted_state122_182_2 + shifted_state122_182_3 + shifted_state122_182_4 + shifted_state122_182_5 + shifted_state122_182_6 + shifted_state122_182_7 + shifted_state122_186_0 + shifted_state122_186_3 + shifted_state122_186_6 + shifted_state122_186_7 + shifted_state122_187_0 + shifted_state122_187_1 + shifted_state122_187_3 + shifted_state122_187_4 + shifted_state122_187_5 + shifted_state122_193_4 + shifted_state122_193_5 + shifted_state122_193_6 + shifted_state122_193_7 + shifted_state122_198_2 + shifted_state122_198_4);
      reservoir_sum_parallel[123] = (shifted_state123_2_0 + shifted_state123_2_1 + shifted_state123_8_4 + shifted_state123_26_0 + shifted_state123_26_1 + shifted_state123_26_5 + shifted_state123_26_6 + shifted_state123_26_7 + shifted_state123_34_0 + shifted_state123_34_1 + shifted_state123_34_3 + shifted_state123_34_4 + shifted_state123_34_5 + shifted_state123_34_6 + shifted_state123_34_7 + shifted_state123_46_0 + shifted_state123_48_0 + shifted_state123_48_1 + shifted_state123_48_4 + shifted_state123_48_6 + shifted_state123_48_7 + shifted_state123_58_6 + shifted_state123_60_0 + shifted_state123_60_1 + shifted_state123_60_3 + shifted_state123_60_4 + shifted_state123_60_6 + shifted_state123_60_7 + shifted_state123_61_2 + shifted_state123_61_3 + shifted_state123_61_5 + shifted_state123_61_6 + shifted_state123_61_7 + shifted_state123_71_3 + shifted_state123_71_5 + shifted_state123_71_6 + shifted_state123_71_7 + shifted_state123_72_0 + shifted_state123_76_4 + shifted_state123_76_6 + shifted_state123_94_4 + shifted_state123_94_5 + shifted_state123_94_7 + shifted_state123_96_4 + shifted_state123_96_5 + shifted_state123_96_6 + shifted_state123_96_7 + shifted_state123_127_1 + shifted_state123_127_2 + shifted_state123_127_3 + shifted_state123_127_4 + shifted_state123_127_5 + shifted_state123_127_6 + shifted_state123_127_7 + shifted_state123_135_0 + shifted_state123_135_1 + shifted_state123_135_5 + shifted_state123_135_6 + shifted_state123_135_7 + shifted_state123_137_3 + shifted_state123_137_6 + shifted_state123_137_7 + shifted_state123_152_0 + shifted_state123_152_1 + shifted_state123_152_2 + shifted_state123_152_3 + shifted_state123_152_4 + shifted_state123_152_5 + shifted_state123_152_6 + shifted_state123_152_7 + shifted_state123_177_0 + shifted_state123_177_1 + shifted_state123_177_2 + shifted_state123_177_4 + shifted_state123_184_0 + shifted_state123_184_3 + shifted_state123_184_4 + shifted_state123_184_5 + shifted_state123_184_6 + shifted_state123_184_7);
      reservoir_sum_parallel[124] = (shifted_state124_0_0 + shifted_state124_0_2 + shifted_state124_0_3 + shifted_state124_0_4 + shifted_state124_0_5 + shifted_state124_0_6 + shifted_state124_0_7 + shifted_state124_21_0 + shifted_state124_21_2 + shifted_state124_21_5 + shifted_state124_21_6 + shifted_state124_21_7 + shifted_state124_38_0 + shifted_state124_38_1 + shifted_state124_38_3 + shifted_state124_38_4 + shifted_state124_38_5 + shifted_state124_38_6 + shifted_state124_38_7 + shifted_state124_53_4 + shifted_state124_55_0 + shifted_state124_55_1 + shifted_state124_55_4 + shifted_state124_55_5 + shifted_state124_55_6 + shifted_state124_55_7 + shifted_state124_57_0 + shifted_state124_57_1 + shifted_state124_57_2 + shifted_state124_57_4 + shifted_state124_57_5 + shifted_state124_57_7 + shifted_state124_71_0 + shifted_state124_71_2 + shifted_state124_71_4 + shifted_state124_71_6 + shifted_state124_71_7 + shifted_state124_76_0 + shifted_state124_76_2 + shifted_state124_76_3 + shifted_state124_76_6 + shifted_state124_76_7 + shifted_state124_80_2 + shifted_state124_80_4 + shifted_state124_100_0 + shifted_state124_100_1 + shifted_state124_100_2 + shifted_state124_100_3 + shifted_state124_100_4 + shifted_state124_100_5 + shifted_state124_100_6 + shifted_state124_100_7 + shifted_state124_109_4 + shifted_state124_109_5 + shifted_state124_109_6 + shifted_state124_109_7 + shifted_state124_114_0 + shifted_state124_114_3 + shifted_state124_114_4 + shifted_state124_119_0 + shifted_state124_119_2 + shifted_state124_119_4 + shifted_state124_119_5 + shifted_state124_119_6 + shifted_state124_119_7 + shifted_state124_136_1 + shifted_state124_136_2 + shifted_state124_136_4 + shifted_state124_142_0 + shifted_state124_142_3 + shifted_state124_142_4 + shifted_state124_142_5 + shifted_state124_142_6 + shifted_state124_142_7 + shifted_state124_151_1 + shifted_state124_151_2 + shifted_state124_151_3 + shifted_state124_151_5 + shifted_state124_160_0 + shifted_state124_160_3 + shifted_state124_160_5 + shifted_state124_160_6 + shifted_state124_160_7 + shifted_state124_162_1 + shifted_state124_162_2 + shifted_state124_162_3 + shifted_state124_185_2 + shifted_state124_185_5 + shifted_state124_185_6 + shifted_state124_185_7 + shifted_state124_186_2 + shifted_state124_186_5 + shifted_state124_186_6 + shifted_state124_186_7 + shifted_state124_189_0 + shifted_state124_189_2 + shifted_state124_189_3 + shifted_state124_189_4 + shifted_state124_189_5 + shifted_state124_189_6 + shifted_state124_189_7 + shifted_state124_196_0 + shifted_state124_196_3 + shifted_state124_196_4 + shifted_state124_198_1 + shifted_state124_198_3);
      reservoir_sum_parallel[125] = (shifted_state125_0_0 + shifted_state125_0_2 + shifted_state125_0_3 + shifted_state125_0_5 + shifted_state125_0_6 + shifted_state125_0_7 + shifted_state125_8_0 + shifted_state125_8_4 + shifted_state125_8_6 + shifted_state125_8_7 + shifted_state125_21_0 + shifted_state125_21_1 + shifted_state125_21_5 + shifted_state125_21_6 + shifted_state125_21_7 + shifted_state125_47_0 + shifted_state125_47_1 + shifted_state125_47_2 + shifted_state125_47_6 + shifted_state125_51_1 + shifted_state125_59_4 + shifted_state125_64_5 + shifted_state125_69_0 + shifted_state125_69_4 + shifted_state125_71_2 + shifted_state125_71_4 + shifted_state125_79_1 + shifted_state125_79_3 + shifted_state125_79_4 + shifted_state125_84_0 + shifted_state125_84_2 + shifted_state125_84_4 + shifted_state125_84_5 + shifted_state125_84_6 + shifted_state125_84_7 + shifted_state125_90_3 + shifted_state125_90_4 + shifted_state125_90_5 + shifted_state125_95_0 + shifted_state125_95_2 + shifted_state125_95_3 + shifted_state125_101_0 + shifted_state125_101_1 + shifted_state125_101_4 + shifted_state125_101_6 + shifted_state125_101_7 + shifted_state125_124_1 + shifted_state125_124_2 + shifted_state125_124_3 + shifted_state125_124_4 + shifted_state125_132_0 + shifted_state125_132_4 + shifted_state125_132_5 + shifted_state125_137_0 + shifted_state125_137_2 + shifted_state125_177_1 + shifted_state125_177_2 + shifted_state125_177_4 + shifted_state125_178_0 + shifted_state125_178_1 + shifted_state125_178_2 + shifted_state125_178_4 + shifted_state125_184_1 + shifted_state125_184_4 + shifted_state125_184_5 + shifted_state125_184_6 + shifted_state125_184_7 + shifted_state125_189_0 + shifted_state125_189_5 + shifted_state125_194_0 + shifted_state125_194_2 + shifted_state125_194_4 + shifted_state125_194_5 + shifted_state125_194_6 + shifted_state125_194_7);
      reservoir_sum_parallel[126] = (shifted_state126_24_0 + shifted_state126_24_2 + shifted_state126_24_3 + shifted_state126_33_0 + shifted_state126_33_2 + shifted_state126_33_3 + shifted_state126_33_5 + shifted_state126_33_6 + shifted_state126_33_7 + shifted_state126_40_2 + shifted_state126_40_3 + shifted_state126_40_5 + shifted_state126_40_6 + shifted_state126_40_7 + shifted_state126_41_0 + shifted_state126_41_3 + shifted_state126_51_0 + shifted_state126_51_3 + shifted_state126_51_4 + shifted_state126_81_0 + shifted_state126_81_1 + shifted_state126_81_2 + shifted_state126_81_4 + shifted_state126_81_6 + shifted_state126_81_7 + shifted_state126_106_0 + shifted_state126_106_1 + shifted_state126_106_2 + shifted_state126_106_3 + shifted_state126_109_1 + shifted_state126_109_5 + shifted_state126_109_6 + shifted_state126_109_7 + shifted_state126_110_1 + shifted_state126_110_2 + shifted_state126_110_4 + shifted_state126_110_5 + shifted_state126_110_6 + shifted_state126_110_7 + shifted_state126_114_0 + shifted_state126_114_3 + shifted_state126_114_4 + shifted_state126_129_1 + shifted_state126_129_2 + shifted_state126_129_5 + shifted_state126_129_6 + shifted_state126_129_7 + shifted_state126_137_0 + shifted_state126_137_1 + shifted_state126_137_3 + shifted_state126_137_4 + shifted_state126_137_6 + shifted_state126_137_7 + shifted_state126_151_2 + shifted_state126_158_1 + shifted_state126_158_3 + shifted_state126_158_4 + shifted_state126_158_5 + shifted_state126_160_0 + shifted_state126_160_3 + shifted_state126_160_4 + shifted_state126_160_5 + shifted_state126_160_6 + shifted_state126_160_7 + shifted_state126_163_5 + shifted_state126_164_0 + shifted_state126_164_1 + shifted_state126_164_2 + shifted_state126_164_4 + shifted_state126_164_5 + shifted_state126_164_6 + shifted_state126_164_7);
      reservoir_sum_parallel[127] = (shifted_state127_8_0 + shifted_state127_8_1 + shifted_state127_8_2 + shifted_state127_8_4 + shifted_state127_17_1 + shifted_state127_17_2 + shifted_state127_17_3 + shifted_state127_17_4 + shifted_state127_17_5 + shifted_state127_17_6 + shifted_state127_17_7 + shifted_state127_26_0 + shifted_state127_26_1 + shifted_state127_26_2 + shifted_state127_26_4 + shifted_state127_42_0 + shifted_state127_42_2 + shifted_state127_42_5 + shifted_state127_42_6 + shifted_state127_42_7 + shifted_state127_51_0 + shifted_state127_51_2 + shifted_state127_51_3 + shifted_state127_51_4 + shifted_state127_51_5 + shifted_state127_54_1 + shifted_state127_54_3 + shifted_state127_104_3 + shifted_state127_165_1 + shifted_state127_165_2 + shifted_state127_165_4 + shifted_state127_165_5 + shifted_state127_168_0 + shifted_state127_168_3 + shifted_state127_168_4 + shifted_state127_168_6 + shifted_state127_168_7 + shifted_state127_174_0 + shifted_state127_174_5 + shifted_state127_174_6 + shifted_state127_174_7);
      reservoir_sum_parallel[128] = (shifted_state128_77_0 + shifted_state128_77_2 + shifted_state128_77_3 + shifted_state128_77_5 + shifted_state128_77_6 + shifted_state128_77_7 + shifted_state128_78_0 + shifted_state128_78_1 + shifted_state128_78_5 + shifted_state128_91_1 + shifted_state128_91_2 + shifted_state128_91_3 + shifted_state128_98_0 + shifted_state128_98_1 + shifted_state128_98_2 + shifted_state128_98_4 + shifted_state128_113_0 + shifted_state128_113_2 + shifted_state128_113_3 + shifted_state128_113_5 + shifted_state128_114_0 + shifted_state128_114_1 + shifted_state128_114_2 + shifted_state128_114_4 + shifted_state128_119_3 + shifted_state128_128_1 + shifted_state128_128_2 + shifted_state128_128_3 + shifted_state128_128_4 + shifted_state128_128_5 + shifted_state128_128_6 + shifted_state128_128_7 + shifted_state128_129_1 + shifted_state128_129_2 + shifted_state128_129_4 + shifted_state128_138_0 + shifted_state128_138_2 + shifted_state128_145_0 + shifted_state128_145_1 + shifted_state128_145_2 + shifted_state128_145_4 + shifted_state128_145_5 + shifted_state128_145_6 + shifted_state128_145_7 + shifted_state128_150_1 + shifted_state128_150_5 + shifted_state128_150_6 + shifted_state128_150_7 + shifted_state128_168_2 + shifted_state128_187_0 + shifted_state128_187_2 + shifted_state128_187_3 + shifted_state128_187_6);
      reservoir_sum_parallel[129] = (shifted_state129_16_0 + shifted_state129_16_1 + shifted_state129_34_0 + shifted_state129_34_1 + shifted_state129_34_3 + shifted_state129_35_0 + shifted_state129_35_2 + shifted_state129_35_5 + shifted_state129_35_7 + shifted_state129_63_0 + shifted_state129_63_1 + shifted_state129_63_3 + shifted_state129_63_4 + shifted_state129_63_5 + shifted_state129_63_6 + shifted_state129_63_7 + shifted_state129_99_2 + shifted_state129_99_3 + shifted_state129_99_4 + shifted_state129_99_6 + shifted_state129_99_7 + shifted_state129_105_0 + shifted_state129_105_1 + shifted_state129_105_3 + shifted_state129_105_5 + shifted_state129_105_6 + shifted_state129_105_7 + shifted_state129_123_0 + shifted_state129_123_3 + shifted_state129_123_5 + shifted_state129_123_6 + shifted_state129_123_7 + shifted_state129_130_1 + shifted_state129_130_2 + shifted_state129_130_4 + shifted_state129_130_5 + shifted_state129_130_6 + shifted_state129_130_7 + shifted_state129_138_3 + shifted_state129_138_4 + shifted_state129_138_5 + shifted_state129_138_6 + shifted_state129_138_7 + shifted_state129_153_0 + shifted_state129_153_1 + shifted_state129_153_2 + shifted_state129_153_4 + shifted_state129_153_5 + shifted_state129_153_6 + shifted_state129_153_7 + shifted_state129_175_2 + shifted_state129_175_3 + shifted_state129_175_5 + shifted_state129_175_6 + shifted_state129_175_7 + shifted_state129_177_0 + shifted_state129_177_2 + shifted_state129_177_3 + shifted_state129_177_4 + shifted_state129_188_0 + shifted_state129_188_3 + shifted_state129_188_4 + shifted_state129_188_5 + shifted_state129_188_6 + shifted_state129_188_7);
      reservoir_sum_parallel[130] = (shifted_state130_23_3 + shifted_state130_24_0 + shifted_state130_24_1 + shifted_state130_24_2 + shifted_state130_24_4 + shifted_state130_24_5 + shifted_state130_24_6 + shifted_state130_24_7 + shifted_state130_37_0 + shifted_state130_37_1 + shifted_state130_37_2 + shifted_state130_37_4 + shifted_state130_38_2 + shifted_state130_50_0 + shifted_state130_50_1 + shifted_state130_50_2 + shifted_state130_50_3 + shifted_state130_50_5 + shifted_state130_50_6 + shifted_state130_50_7 + shifted_state130_63_0 + shifted_state130_63_1 + shifted_state130_63_2 + shifted_state130_63_3 + shifted_state130_63_4 + shifted_state130_63_5 + shifted_state130_63_6 + shifted_state130_63_7 + shifted_state130_78_1 + shifted_state130_78_2 + shifted_state130_78_3 + shifted_state130_78_4 + shifted_state130_78_6 + shifted_state130_78_7 + shifted_state130_80_3 + shifted_state130_80_4 + shifted_state130_80_6 + shifted_state130_80_7 + shifted_state130_85_2 + shifted_state130_85_3 + shifted_state130_97_1 + shifted_state130_97_2 + shifted_state130_104_4 + shifted_state130_104_5 + shifted_state130_104_6 + shifted_state130_104_7 + shifted_state130_116_3 + shifted_state130_116_5 + shifted_state130_116_6 + shifted_state130_116_7 + shifted_state130_118_1 + shifted_state130_118_2 + shifted_state130_118_3 + shifted_state130_146_0 + shifted_state130_146_2 + shifted_state130_146_4 + shifted_state130_146_5 + shifted_state130_146_6 + shifted_state130_146_7 + shifted_state130_152_0 + shifted_state130_152_1 + shifted_state130_164_0 + shifted_state130_164_4 + shifted_state130_164_5 + shifted_state130_164_6 + shifted_state130_164_7 + shifted_state130_167_0 + shifted_state130_169_0 + shifted_state130_169_4 + shifted_state130_177_5 + shifted_state130_177_6 + shifted_state130_177_7 + shifted_state130_181_0 + shifted_state130_181_1 + shifted_state130_181_3 + shifted_state130_181_6 + shifted_state130_181_7 + shifted_state130_191_0 + shifted_state130_191_1 + shifted_state130_191_2 + shifted_state130_191_3 + shifted_state130_191_4 + shifted_state130_192_0 + shifted_state130_192_1 + shifted_state130_192_4 + shifted_state130_192_6 + shifted_state130_192_7);
      reservoir_sum_parallel[131] = (shifted_state131_13_1 + shifted_state131_19_2 + shifted_state131_19_3 + shifted_state131_20_0 + shifted_state131_20_5 + shifted_state131_20_6 + shifted_state131_20_7 + shifted_state131_25_1 + shifted_state131_25_2 + shifted_state131_25_5 + shifted_state131_25_6 + shifted_state131_25_7 + shifted_state131_28_0 + shifted_state131_28_1 + shifted_state131_28_3 + shifted_state131_28_5 + shifted_state131_31_1 + shifted_state131_31_2 + shifted_state131_31_3 + shifted_state131_50_0 + shifted_state131_50_2 + shifted_state131_50_3 + shifted_state131_56_3 + shifted_state131_56_4 + shifted_state131_56_5 + shifted_state131_56_6 + shifted_state131_56_7 + shifted_state131_71_0 + shifted_state131_71_1 + shifted_state131_71_2 + shifted_state131_71_5 + shifted_state131_71_6 + shifted_state131_71_7 + shifted_state131_72_2 + shifted_state131_72_3 + shifted_state131_72_5 + shifted_state131_72_6 + shifted_state131_72_7 + shifted_state131_74_2 + shifted_state131_74_4 + shifted_state131_74_6 + shifted_state131_74_7 + shifted_state131_76_0 + shifted_state131_76_2 + shifted_state131_76_3 + shifted_state131_99_0 + shifted_state131_99_5 + shifted_state131_99_6 + shifted_state131_99_7 + shifted_state131_106_0 + shifted_state131_106_1 + shifted_state131_106_4 + shifted_state131_118_0 + shifted_state131_118_1 + shifted_state131_118_2 + shifted_state131_118_3 + shifted_state131_118_4 + shifted_state131_118_6 + shifted_state131_118_7 + shifted_state131_121_0 + shifted_state131_121_3 + shifted_state131_121_5 + shifted_state131_121_6 + shifted_state131_121_7 + shifted_state131_127_2 + shifted_state131_127_5 + shifted_state131_133_0 + shifted_state131_133_3 + shifted_state131_133_4 + shifted_state131_134_1 + shifted_state131_134_2 + shifted_state131_134_3 + shifted_state131_134_6 + shifted_state131_155_1 + shifted_state131_155_4 + shifted_state131_174_2 + shifted_state131_174_3 + shifted_state131_175_1 + shifted_state131_175_2 + shifted_state131_175_3 + shifted_state131_175_4);
      reservoir_sum_parallel[132] = (shifted_state132_4_0 + shifted_state132_4_1 + shifted_state132_4_2 + shifted_state132_4_3 + shifted_state132_4_4 + shifted_state132_4_5 + shifted_state132_4_6 + shifted_state132_4_7 + shifted_state132_16_1 + shifted_state132_16_4 + shifted_state132_16_5 + shifted_state132_16_6 + shifted_state132_16_7 + shifted_state132_19_0 + shifted_state132_19_2 + shifted_state132_19_4 + shifted_state132_19_5 + shifted_state132_19_6 + shifted_state132_19_7 + shifted_state132_32_1 + shifted_state132_32_4 + shifted_state132_33_0 + shifted_state132_33_5 + shifted_state132_35_1 + shifted_state132_35_2 + shifted_state132_35_3 + shifted_state132_35_4 + shifted_state132_35_5 + shifted_state132_35_6 + shifted_state132_35_7 + shifted_state132_48_1 + shifted_state132_48_4 + shifted_state132_48_6 + shifted_state132_60_0 + shifted_state132_60_2 + shifted_state132_60_3 + shifted_state132_60_4 + shifted_state132_60_5 + shifted_state132_60_6 + shifted_state132_60_7 + shifted_state132_65_0 + shifted_state132_65_5 + shifted_state132_67_5 + shifted_state132_102_0 + shifted_state132_102_2 + shifted_state132_102_3 + shifted_state132_102_4 + shifted_state132_122_1 + shifted_state132_122_3 + shifted_state132_122_5 + shifted_state132_126_3 + shifted_state132_126_4 + shifted_state132_126_5 + shifted_state132_126_6 + shifted_state132_126_7 + shifted_state132_132_1 + shifted_state132_132_5 + shifted_state132_138_0 + shifted_state132_138_3 + shifted_state132_138_5 + shifted_state132_138_6 + shifted_state132_138_7 + shifted_state132_150_0 + shifted_state132_150_1 + shifted_state132_169_3);
      reservoir_sum_parallel[133] = (shifted_state133_5_0 + shifted_state133_5_5 + shifted_state133_38_1 + shifted_state133_38_2 + shifted_state133_38_3 + shifted_state133_38_4 + shifted_state133_40_0 + shifted_state133_40_1 + shifted_state133_40_2 + shifted_state133_40_5 + shifted_state133_40_7 + shifted_state133_51_1 + shifted_state133_51_2 + shifted_state133_55_3 + shifted_state133_55_5 + shifted_state133_55_6 + shifted_state133_55_7 + shifted_state133_66_3 + shifted_state133_68_0 + shifted_state133_68_1 + shifted_state133_68_2 + shifted_state133_68_4 + shifted_state133_68_5 + shifted_state133_68_6 + shifted_state133_68_7 + shifted_state133_80_0 + shifted_state133_80_1 + shifted_state133_80_4 + shifted_state133_80_5 + shifted_state133_84_0 + shifted_state133_84_2 + shifted_state133_84_4 + shifted_state133_84_6 + shifted_state133_84_7 + shifted_state133_88_0 + shifted_state133_88_1 + shifted_state133_88_2 + shifted_state133_88_3 + shifted_state133_88_4 + shifted_state133_92_0 + shifted_state133_92_3 + shifted_state133_92_5 + shifted_state133_111_0 + shifted_state133_111_1 + shifted_state133_111_2 + shifted_state133_111_3 + shifted_state133_111_4 + shifted_state133_139_5 + shifted_state133_156_0 + shifted_state133_156_1 + shifted_state133_156_2 + shifted_state133_156_3 + shifted_state133_156_4 + shifted_state133_167_0 + shifted_state133_167_3 + shifted_state133_167_5 + shifted_state133_168_0 + shifted_state133_168_1 + shifted_state133_168_2 + shifted_state133_168_3 + shifted_state133_168_4 + shifted_state133_168_6 + shifted_state133_175_1 + shifted_state133_175_3 + shifted_state133_175_4 + shifted_state133_175_5 + shifted_state133_176_3 + shifted_state133_176_5 + shifted_state133_176_6 + shifted_state133_176_7 + shifted_state133_190_0 + shifted_state133_190_1 + shifted_state133_190_2 + shifted_state133_190_3 + shifted_state133_190_4 + shifted_state133_190_5 + shifted_state133_190_6 + shifted_state133_190_7 + shifted_state133_194_5 + shifted_state133_199_0 + shifted_state133_199_1 + shifted_state133_199_3);
      reservoir_sum_parallel[134] = (shifted_state134_9_1 + shifted_state134_9_4 + shifted_state134_9_5 + shifted_state134_9_6 + shifted_state134_9_7 + shifted_state134_15_1 + shifted_state134_15_2 + shifted_state134_15_4 + shifted_state134_15_5 + shifted_state134_15_6 + shifted_state134_15_7 + shifted_state134_24_1 + shifted_state134_24_4 + shifted_state134_24_5 + shifted_state134_24_6 + shifted_state134_24_7 + shifted_state134_25_0 + shifted_state134_25_2 + shifted_state134_25_3 + shifted_state134_25_4 + shifted_state134_25_6 + shifted_state134_25_7 + shifted_state134_39_1 + shifted_state134_39_2 + shifted_state134_39_3 + shifted_state134_54_1 + shifted_state134_54_5 + shifted_state134_70_4 + shifted_state134_88_1 + shifted_state134_88_5 + shifted_state134_88_6 + shifted_state134_88_7 + shifted_state134_89_0 + shifted_state134_89_2 + shifted_state134_89_3 + shifted_state134_89_4 + shifted_state134_89_6 + shifted_state134_89_7 + shifted_state134_94_0 + shifted_state134_94_1 + shifted_state134_94_2 + shifted_state134_94_4 + shifted_state134_94_6 + shifted_state134_94_7 + shifted_state134_100_0 + shifted_state134_100_1 + shifted_state134_100_2 + shifted_state134_103_5 + shifted_state134_103_6 + shifted_state134_103_7 + shifted_state134_108_0 + shifted_state134_108_1 + shifted_state134_108_2 + shifted_state134_108_5 + shifted_state134_134_1 + shifted_state134_134_2 + shifted_state134_134_3 + shifted_state134_134_5 + shifted_state134_134_6 + shifted_state134_134_7 + shifted_state134_164_1 + shifted_state134_164_3 + shifted_state134_166_0 + shifted_state134_166_2 + shifted_state134_166_3 + shifted_state134_185_1 + shifted_state134_185_3 + shifted_state134_194_0 + shifted_state134_194_1 + shifted_state134_194_2);
      reservoir_sum_parallel[135] = (shifted_state135_23_0 + shifted_state135_23_2 + shifted_state135_23_3 + shifted_state135_23_4 + shifted_state135_25_0 + shifted_state135_25_2 + shifted_state135_46_0 + shifted_state135_46_4 + shifted_state135_46_5 + shifted_state135_46_6 + shifted_state135_46_7 + shifted_state135_65_0 + shifted_state135_65_1 + shifted_state135_65_2 + shifted_state135_65_3 + shifted_state135_65_4 + shifted_state135_78_2 + shifted_state135_78_3 + shifted_state135_78_5 + shifted_state135_78_6 + shifted_state135_78_7 + shifted_state135_81_2 + shifted_state135_81_3 + shifted_state135_84_1 + shifted_state135_91_1 + shifted_state135_91_2 + shifted_state135_91_5 + shifted_state135_112_0 + shifted_state135_112_1 + shifted_state135_112_4 + shifted_state135_130_1 + shifted_state135_130_2 + shifted_state135_130_5 + shifted_state135_133_1 + shifted_state135_133_2 + shifted_state135_133_5 + shifted_state135_133_6 + shifted_state135_133_7 + shifted_state135_142_0 + shifted_state135_142_3 + shifted_state135_142_4 + shifted_state135_142_5 + shifted_state135_142_6 + shifted_state135_142_7 + shifted_state135_144_1 + shifted_state135_144_4 + shifted_state135_144_5 + shifted_state135_144_6 + shifted_state135_144_7 + shifted_state135_161_1 + shifted_state135_161_3 + shifted_state135_161_4 + shifted_state135_161_6 + shifted_state135_161_7 + shifted_state135_164_2 + shifted_state135_164_5 + shifted_state135_168_0 + shifted_state135_168_1 + shifted_state135_168_3 + shifted_state135_168_5 + shifted_state135_168_6 + shifted_state135_168_7 + shifted_state135_182_0 + shifted_state135_182_1 + shifted_state135_182_4 + shifted_state135_190_1 + shifted_state135_190_2 + shifted_state135_190_4 + shifted_state135_190_5 + shifted_state135_190_6 + shifted_state135_190_7 + shifted_state135_191_1 + shifted_state135_191_3 + shifted_state135_191_5 + shifted_state135_191_6 + shifted_state135_191_7);
      reservoir_sum_parallel[136] = (shifted_state136_14_1 + shifted_state136_14_4 + shifted_state136_14_5 + shifted_state136_14_6 + shifted_state136_14_7 + shifted_state136_18_1 + shifted_state136_18_2 + shifted_state136_18_4 + shifted_state136_18_5 + shifted_state136_18_6 + shifted_state136_18_7 + shifted_state136_25_1 + shifted_state136_25_2 + shifted_state136_25_3 + shifted_state136_25_4 + shifted_state136_25_5 + shifted_state136_25_6 + shifted_state136_25_7 + shifted_state136_31_2 + shifted_state136_31_3 + shifted_state136_31_5 + shifted_state136_31_6 + shifted_state136_31_7 + shifted_state136_33_0 + shifted_state136_33_1 + shifted_state136_33_2 + shifted_state136_33_3 + shifted_state136_33_4 + shifted_state136_33_5 + shifted_state136_33_6 + shifted_state136_33_7 + shifted_state136_37_1 + shifted_state136_37_3 + shifted_state136_37_4 + shifted_state136_37_6 + shifted_state136_37_7 + shifted_state136_41_0 + shifted_state136_41_1 + shifted_state136_41_2 + shifted_state136_41_5 + shifted_state136_41_6 + shifted_state136_41_7 + shifted_state136_43_0 + shifted_state136_43_2 + shifted_state136_43_5 + shifted_state136_53_0 + shifted_state136_53_1 + shifted_state136_53_2 + shifted_state136_53_3 + shifted_state136_53_4 + shifted_state136_53_5 + shifted_state136_53_6 + shifted_state136_53_7 + shifted_state136_81_1 + shifted_state136_81_3 + shifted_state136_81_4 + shifted_state136_81_5 + shifted_state136_81_6 + shifted_state136_81_7 + shifted_state136_82_0 + shifted_state136_82_1 + shifted_state136_82_4 + shifted_state136_82_6 + shifted_state136_85_0 + shifted_state136_85_1 + shifted_state136_85_5 + shifted_state136_85_6 + shifted_state136_85_7 + shifted_state136_87_0 + shifted_state136_87_2 + shifted_state136_87_4 + shifted_state136_106_0 + shifted_state136_106_1 + shifted_state136_106_2 + shifted_state136_106_4 + shifted_state136_106_6 + shifted_state136_106_7 + shifted_state136_120_0 + shifted_state136_120_1 + shifted_state136_120_3 + shifted_state136_120_4 + shifted_state136_120_5 + shifted_state136_129_2 + shifted_state136_129_4 + shifted_state136_129_5 + shifted_state136_130_0 + shifted_state136_130_1 + shifted_state136_130_5 + shifted_state136_136_0 + shifted_state136_136_1 + shifted_state136_136_3 + shifted_state136_136_5 + shifted_state136_139_1 + shifted_state136_139_5 + shifted_state136_139_6 + shifted_state136_139_7 + shifted_state136_141_0 + shifted_state136_141_1 + shifted_state136_141_2 + shifted_state136_141_4 + shifted_state136_141_5 + shifted_state136_180_0 + shifted_state136_180_1 + shifted_state136_180_3 + shifted_state136_191_4 + shifted_state136_191_5 + shifted_state136_191_7);
      reservoir_sum_parallel[137] = (shifted_state137_8_0 + shifted_state137_8_5 + shifted_state137_9_5 + shifted_state137_9_6 + shifted_state137_9_7 + shifted_state137_23_4 + shifted_state137_23_5 + shifted_state137_23_6 + shifted_state137_23_7 + shifted_state137_28_2 + shifted_state137_28_3 + shifted_state137_40_1 + shifted_state137_40_3 + shifted_state137_40_5 + shifted_state137_40_6 + shifted_state137_40_7 + shifted_state137_51_1 + shifted_state137_51_4 + shifted_state137_51_5 + shifted_state137_51_6 + shifted_state137_51_7 + shifted_state137_52_1 + shifted_state137_52_4 + shifted_state137_54_0 + shifted_state137_54_1 + shifted_state137_54_5 + shifted_state137_63_2 + shifted_state137_63_3 + shifted_state137_66_0 + shifted_state137_66_2 + shifted_state137_66_4 + shifted_state137_66_6 + shifted_state137_66_7 + shifted_state137_78_0 + shifted_state137_78_2 + shifted_state137_92_0 + shifted_state137_92_3 + shifted_state137_92_4 + shifted_state137_92_5 + shifted_state137_92_6 + shifted_state137_92_7 + shifted_state137_101_0 + shifted_state137_101_5 + shifted_state137_101_6 + shifted_state137_101_7 + shifted_state137_103_0 + shifted_state137_103_3 + shifted_state137_103_5 + shifted_state137_106_3 + shifted_state137_106_4 + shifted_state137_106_5 + shifted_state137_106_6 + shifted_state137_106_7 + shifted_state137_112_0 + shifted_state137_112_1 + shifted_state137_112_5 + shifted_state137_114_3 + shifted_state137_114_4 + shifted_state137_114_5 + shifted_state137_114_6 + shifted_state137_114_7 + shifted_state137_115_0 + shifted_state137_115_4 + shifted_state137_115_6 + shifted_state137_115_7 + shifted_state137_141_0 + shifted_state137_141_1 + shifted_state137_141_2 + shifted_state137_141_3 + shifted_state137_141_4 + shifted_state137_141_6 + shifted_state137_141_7 + shifted_state137_158_4 + shifted_state137_158_5 + shifted_state137_158_7 + shifted_state137_175_1 + shifted_state137_175_2 + shifted_state137_175_3 + shifted_state137_175_4 + shifted_state137_175_6 + shifted_state137_175_7 + shifted_state137_182_1 + shifted_state137_182_2 + shifted_state137_182_3 + shifted_state137_188_0 + shifted_state137_188_1 + shifted_state137_188_2 + shifted_state137_188_3 + shifted_state137_188_5 + shifted_state137_188_6 + shifted_state137_188_7);
      reservoir_sum_parallel[138] = (shifted_state138_19_2 + shifted_state138_19_3 + shifted_state138_20_5 + shifted_state138_20_6 + shifted_state138_20_7 + shifted_state138_26_0 + shifted_state138_26_3 + shifted_state138_26_5 + shifted_state138_26_6 + shifted_state138_26_7 + shifted_state138_28_3 + shifted_state138_54_0 + shifted_state138_54_2 + shifted_state138_54_5 + shifted_state138_72_0 + shifted_state138_72_1 + shifted_state138_72_3 + shifted_state138_72_4 + shifted_state138_72_5 + shifted_state138_81_0 + shifted_state138_81_1 + shifted_state138_81_2 + shifted_state138_81_3 + shifted_state138_81_4 + shifted_state138_81_5 + shifted_state138_81_6 + shifted_state138_81_7 + shifted_state138_85_0 + shifted_state138_85_1 + shifted_state138_85_5 + shifted_state138_85_6 + shifted_state138_85_7 + shifted_state138_94_0 + shifted_state138_94_1 + shifted_state138_94_2 + shifted_state138_94_3 + shifted_state138_104_2 + shifted_state138_104_4 + shifted_state138_104_5 + shifted_state138_104_7 + shifted_state138_107_1 + shifted_state138_107_2 + shifted_state138_107_3 + shifted_state138_125_0 + shifted_state138_125_4 + shifted_state138_140_1 + shifted_state138_140_2 + shifted_state138_140_3 + shifted_state138_140_4 + shifted_state138_144_1 + shifted_state138_144_2 + shifted_state138_144_5 + shifted_state138_144_6 + shifted_state138_144_7 + shifted_state138_149_3 + shifted_state138_149_4 + shifted_state138_149_5 + shifted_state138_149_6 + shifted_state138_149_7 + shifted_state138_150_0 + shifted_state138_150_3 + shifted_state138_150_4 + shifted_state138_158_1 + shifted_state138_158_2 + shifted_state138_158_3 + shifted_state138_158_4 + shifted_state138_163_1 + shifted_state138_163_3 + shifted_state138_163_4 + shifted_state138_163_5 + shifted_state138_163_6 + shifted_state138_163_7 + shifted_state138_177_2 + shifted_state138_177_3 + shifted_state138_177_5 + shifted_state138_177_6 + shifted_state138_177_7 + shifted_state138_183_1 + shifted_state138_183_3 + shifted_state138_183_5 + shifted_state138_183_6 + shifted_state138_183_7 + shifted_state138_192_0 + shifted_state138_192_1 + shifted_state138_192_2 + shifted_state138_192_3 + shifted_state138_192_4 + shifted_state138_193_0 + shifted_state138_193_3);
      reservoir_sum_parallel[139] = (shifted_state139_19_0 + shifted_state139_19_4 + shifted_state139_19_5 + shifted_state139_46_0 + shifted_state139_46_3 + shifted_state139_49_0 + shifted_state139_49_2 + shifted_state139_49_4 + shifted_state139_49_5 + shifted_state139_49_6 + shifted_state139_49_7 + shifted_state139_56_0 + shifted_state139_56_3 + shifted_state139_56_4 + shifted_state139_56_6 + shifted_state139_56_7 + shifted_state139_61_1 + shifted_state139_61_2 + shifted_state139_61_3 + shifted_state139_61_5 + shifted_state139_78_0 + shifted_state139_78_2 + shifted_state139_78_3 + shifted_state139_78_5 + shifted_state139_78_6 + shifted_state139_78_7 + shifted_state139_89_1 + shifted_state139_89_2 + shifted_state139_89_5 + shifted_state139_89_6 + shifted_state139_89_7 + shifted_state139_97_0 + shifted_state139_97_3 + shifted_state139_97_5 + shifted_state139_97_6 + shifted_state139_97_7 + shifted_state139_141_0 + shifted_state139_141_1 + shifted_state139_141_2 + shifted_state139_141_4 + shifted_state139_141_5 + shifted_state139_151_0 + shifted_state139_151_1 + shifted_state139_151_3 + shifted_state139_151_4 + shifted_state139_151_5 + shifted_state139_157_2 + shifted_state139_157_3 + shifted_state139_157_4 + shifted_state139_157_6 + shifted_state139_157_7 + shifted_state139_178_3 + shifted_state139_178_5 + shifted_state139_185_0 + shifted_state139_185_2 + shifted_state139_185_4 + shifted_state139_191_0 + shifted_state139_191_4);
      reservoir_sum_parallel[140] = (shifted_state140_4_3 + shifted_state140_4_5 + shifted_state140_21_2 + shifted_state140_21_4 + shifted_state140_21_5 + shifted_state140_27_2 + shifted_state140_27_4 + shifted_state140_38_0 + shifted_state140_38_2 + shifted_state140_38_3 + shifted_state140_38_6 + shifted_state140_38_7 + shifted_state140_43_0 + shifted_state140_43_2 + shifted_state140_44_1 + shifted_state140_44_2 + shifted_state140_44_3 + shifted_state140_44_4 + shifted_state140_64_1 + shifted_state140_64_2 + shifted_state140_64_3 + shifted_state140_83_0 + shifted_state140_83_1 + shifted_state140_83_2 + shifted_state140_83_5 + shifted_state140_83_6 + shifted_state140_83_7 + shifted_state140_94_3 + shifted_state140_94_4 + shifted_state140_94_6 + shifted_state140_94_7 + shifted_state140_104_0 + shifted_state140_121_0 + shifted_state140_121_2 + shifted_state140_121_6 + shifted_state140_121_7 + shifted_state140_129_0 + shifted_state140_129_2 + shifted_state140_129_4 + shifted_state140_133_0 + shifted_state140_133_2 + shifted_state140_133_4 + shifted_state140_138_1 + shifted_state140_138_2 + shifted_state140_138_3 + shifted_state140_138_5 + shifted_state140_138_6 + shifted_state140_138_7 + shifted_state140_152_0 + shifted_state140_152_2 + shifted_state140_152_4 + shifted_state140_155_1 + shifted_state140_155_2 + shifted_state140_155_3 + shifted_state140_155_4 + shifted_state140_155_5 + shifted_state140_155_6 + shifted_state140_155_7 + shifted_state140_165_0 + shifted_state140_165_1 + shifted_state140_165_3 + shifted_state140_165_6 + shifted_state140_165_7 + shifted_state140_174_0 + shifted_state140_174_4 + shifted_state140_182_0 + shifted_state140_182_1 + shifted_state140_182_2 + shifted_state140_182_5 + shifted_state140_183_3 + shifted_state140_183_4);
      reservoir_sum_parallel[141] = (shifted_state141_7_1 + shifted_state141_7_2 + shifted_state141_7_5 + shifted_state141_7_6 + shifted_state141_7_7 + shifted_state141_11_1 + shifted_state141_11_2 + shifted_state141_11_3 + shifted_state141_13_0 + shifted_state141_13_3 + shifted_state141_16_4 + shifted_state141_32_1 + shifted_state141_32_2 + shifted_state141_32_3 + shifted_state141_32_5 + shifted_state141_35_2 + shifted_state141_35_3 + shifted_state141_37_2 + shifted_state141_37_5 + shifted_state141_37_6 + shifted_state141_37_7 + shifted_state141_41_0 + shifted_state141_41_3 + shifted_state141_41_4 + shifted_state141_41_5 + shifted_state141_46_0 + shifted_state141_46_1 + shifted_state141_46_3 + shifted_state141_46_5 + shifted_state141_53_0 + shifted_state141_53_2 + shifted_state141_53_5 + shifted_state141_53_6 + shifted_state141_53_7 + shifted_state141_65_6 + shifted_state141_65_7 + shifted_state141_75_0 + shifted_state141_85_0 + shifted_state141_85_2 + shifted_state141_85_3 + shifted_state141_97_3 + shifted_state141_97_5 + shifted_state141_97_6 + shifted_state141_97_7 + shifted_state141_109_0 + shifted_state141_109_1 + shifted_state141_109_2 + shifted_state141_109_4 + shifted_state141_109_6 + shifted_state141_109_7 + shifted_state141_112_0 + shifted_state141_112_4 + shifted_state141_112_6 + shifted_state141_112_7 + shifted_state141_125_0 + shifted_state141_125_1 + shifted_state141_125_3 + shifted_state141_127_0 + shifted_state141_127_1 + shifted_state141_127_3 + shifted_state141_127_5 + shifted_state141_131_0 + shifted_state141_131_1 + shifted_state141_131_2 + shifted_state141_131_3 + shifted_state141_131_5 + shifted_state141_148_4 + shifted_state141_150_0 + shifted_state141_150_1 + shifted_state141_150_3 + shifted_state141_150_6 + shifted_state141_150_7 + shifted_state141_151_0 + shifted_state141_151_1 + shifted_state141_151_3 + shifted_state141_152_1 + shifted_state141_160_0 + shifted_state141_160_2 + shifted_state141_160_4 + shifted_state141_160_6 + shifted_state141_160_7 + shifted_state141_171_0 + shifted_state141_171_2 + shifted_state141_171_4 + shifted_state141_171_6 + shifted_state141_171_7 + shifted_state141_184_0 + shifted_state141_184_1 + shifted_state141_184_3 + shifted_state141_184_4 + shifted_state141_184_6 + shifted_state141_184_7 + shifted_state141_189_0 + shifted_state141_189_4 + shifted_state141_192_0 + shifted_state141_192_3 + shifted_state141_192_5 + shifted_state141_197_0 + shifted_state141_197_5 + shifted_state141_197_6 + shifted_state141_197_7);
      reservoir_sum_parallel[142] = (shifted_state142_5_1 + shifted_state142_5_3 + shifted_state142_5_4 + shifted_state142_44_0 + shifted_state142_44_2 + shifted_state142_44_3 + shifted_state142_44_5 + shifted_state142_44_6 + shifted_state142_44_7 + shifted_state142_46_1 + shifted_state142_46_2 + shifted_state142_46_4 + shifted_state142_46_5 + shifted_state142_46_6 + shifted_state142_46_7 + shifted_state142_49_2 + shifted_state142_49_3 + shifted_state142_49_4 + shifted_state142_49_5 + shifted_state142_49_6 + shifted_state142_49_7 + shifted_state142_51_0 + shifted_state142_51_1 + shifted_state142_51_3 + shifted_state142_53_0 + shifted_state142_53_1 + shifted_state142_53_2 + shifted_state142_53_6 + shifted_state142_59_0 + shifted_state142_65_0 + shifted_state142_65_3 + shifted_state142_65_4 + shifted_state142_71_0 + shifted_state142_71_1 + shifted_state142_71_2 + shifted_state142_71_6 + shifted_state142_71_7 + shifted_state142_73_1 + shifted_state142_73_2 + shifted_state142_73_3 + shifted_state142_73_4 + shifted_state142_73_6 + shifted_state142_73_7 + shifted_state142_76_0 + shifted_state142_76_2 + shifted_state142_81_1 + shifted_state142_81_3 + shifted_state142_84_0 + shifted_state142_84_1 + shifted_state142_84_3 + shifted_state142_84_4 + shifted_state142_99_1 + shifted_state142_99_2 + shifted_state142_99_4 + shifted_state142_100_0 + shifted_state142_100_4 + shifted_state142_100_6 + shifted_state142_100_7 + shifted_state142_113_0 + shifted_state142_113_1 + shifted_state142_113_2 + shifted_state142_113_3 + shifted_state142_113_5 + shifted_state142_124_0 + shifted_state142_124_1 + shifted_state142_124_4 + shifted_state142_125_1 + shifted_state142_125_4 + shifted_state142_125_5 + shifted_state142_131_1 + shifted_state142_131_3 + shifted_state142_131_4 + shifted_state142_131_6 + shifted_state142_131_7 + shifted_state142_138_1 + shifted_state142_138_3 + shifted_state142_138_4 + shifted_state142_138_5 + shifted_state142_144_1 + shifted_state142_144_2 + shifted_state142_156_1 + shifted_state142_156_2 + shifted_state142_156_5 + shifted_state142_179_1 + shifted_state142_179_3 + shifted_state142_191_0 + shifted_state142_191_1 + shifted_state142_191_2 + shifted_state142_191_4 + shifted_state142_193_0 + shifted_state142_193_1 + shifted_state142_193_2 + shifted_state142_193_3 + shifted_state142_193_4 + shifted_state142_193_5 + shifted_state142_193_6 + shifted_state142_193_7 + shifted_state142_196_3 + shifted_state142_196_5);
      reservoir_sum_parallel[143] = (shifted_state143_0_0 + shifted_state143_0_1 + shifted_state143_0_2 + shifted_state143_0_4 + shifted_state143_9_1 + shifted_state143_9_2 + shifted_state143_9_3 + shifted_state143_18_1 + shifted_state143_18_2 + shifted_state143_18_5 + shifted_state143_18_6 + shifted_state143_18_7 + shifted_state143_20_0 + shifted_state143_20_2 + shifted_state143_20_3 + shifted_state143_20_4 + shifted_state143_30_2 + shifted_state143_32_0 + shifted_state143_32_1 + shifted_state143_32_2 + shifted_state143_32_3 + shifted_state143_32_4 + shifted_state143_32_5 + shifted_state143_32_6 + shifted_state143_32_7 + shifted_state143_33_0 + shifted_state143_33_1 + shifted_state143_33_3 + shifted_state143_33_4 + shifted_state143_47_3 + shifted_state143_54_1 + shifted_state143_54_2 + shifted_state143_54_5 + shifted_state143_58_0 + shifted_state143_58_1 + shifted_state143_58_3 + shifted_state143_58_5 + shifted_state143_58_6 + shifted_state143_58_7 + shifted_state143_83_1 + shifted_state143_83_3 + shifted_state143_83_4 + shifted_state143_89_1 + shifted_state143_89_3 + shifted_state143_89_6 + shifted_state143_89_7 + shifted_state143_103_0 + shifted_state143_103_6 + shifted_state143_103_7 + shifted_state143_113_0 + shifted_state143_113_1 + shifted_state143_113_2 + shifted_state143_113_3 + shifted_state143_113_4 + shifted_state143_113_5 + shifted_state143_113_6 + shifted_state143_113_7 + shifted_state143_130_0 + shifted_state143_130_1 + shifted_state143_130_3 + shifted_state143_130_6 + shifted_state143_130_7 + shifted_state143_134_2 + shifted_state143_134_5 + shifted_state143_169_0 + shifted_state143_169_1 + shifted_state143_169_4 + shifted_state143_169_6 + shifted_state143_169_7 + shifted_state143_183_3 + shifted_state143_183_4 + shifted_state143_183_6 + shifted_state143_183_7 + shifted_state143_187_1 + shifted_state143_187_6 + shifted_state143_187_7 + shifted_state143_192_0 + shifted_state143_192_3);
      reservoir_sum_parallel[144] = (shifted_state144_14_2 + shifted_state144_14_3 + shifted_state144_14_4 + shifted_state144_14_5 + shifted_state144_14_6 + shifted_state144_14_7 + shifted_state144_15_0 + shifted_state144_15_2 + shifted_state144_16_2 + shifted_state144_44_0 + shifted_state144_44_3 + shifted_state144_44_6 + shifted_state144_44_7 + shifted_state144_49_1 + shifted_state144_49_5 + shifted_state144_51_1 + shifted_state144_51_2 + shifted_state144_51_3 + shifted_state144_51_4 + shifted_state144_51_5 + shifted_state144_51_6 + shifted_state144_51_7 + shifted_state144_84_1 + shifted_state144_84_3 + shifted_state144_84_4 + shifted_state144_100_0 + shifted_state144_100_1 + shifted_state144_100_2 + shifted_state144_100_4 + shifted_state144_100_5 + shifted_state144_109_0 + shifted_state144_109_1 + shifted_state144_109_2 + shifted_state144_109_6 + shifted_state144_125_1 + shifted_state144_125_3 + shifted_state144_125_6 + shifted_state144_125_7 + shifted_state144_128_0 + shifted_state144_128_1 + shifted_state144_128_2 + shifted_state144_134_4 + shifted_state144_135_0 + shifted_state144_135_1 + shifted_state144_135_2 + shifted_state144_135_3 + shifted_state144_135_5 + shifted_state144_139_2 + shifted_state144_139_3 + shifted_state144_139_4 + shifted_state144_142_0 + shifted_state144_142_1 + shifted_state144_142_2 + shifted_state144_142_3 + shifted_state144_142_5 + shifted_state144_142_6 + shifted_state144_142_7 + shifted_state144_166_0 + shifted_state144_166_2 + shifted_state144_166_3 + shifted_state144_166_5 + shifted_state144_166_6 + shifted_state144_166_7 + shifted_state144_181_0 + shifted_state144_181_1 + shifted_state144_181_3 + shifted_state144_184_0 + shifted_state144_184_3 + shifted_state144_184_5 + shifted_state144_184_6 + shifted_state144_184_7);
      reservoir_sum_parallel[145] = (shifted_state145_13_0 + shifted_state145_22_0 + shifted_state145_22_3 + shifted_state145_22_4 + shifted_state145_24_0 + shifted_state145_24_2 + shifted_state145_24_4 + shifted_state145_31_0 + shifted_state145_31_2 + shifted_state145_31_3 + shifted_state145_31_6 + shifted_state145_31_7 + shifted_state145_43_0 + shifted_state145_43_3 + shifted_state145_43_4 + shifted_state145_43_5 + shifted_state145_43_7 + shifted_state145_45_0 + shifted_state145_45_3 + shifted_state145_45_4 + shifted_state145_49_4 + shifted_state145_51_1 + shifted_state145_51_3 + shifted_state145_68_1 + shifted_state145_68_2 + shifted_state145_68_4 + shifted_state145_68_5 + shifted_state145_68_7 + shifted_state145_74_1 + shifted_state145_74_2 + shifted_state145_74_5 + shifted_state145_74_6 + shifted_state145_74_7 + shifted_state145_97_4 + shifted_state145_97_5 + shifted_state145_97_6 + shifted_state145_97_7 + shifted_state145_109_0 + shifted_state145_109_1 + shifted_state145_109_3 + shifted_state145_109_5 + shifted_state145_116_0 + shifted_state145_116_2 + shifted_state145_116_3 + shifted_state145_116_4 + shifted_state145_126_2 + shifted_state145_126_4 + shifted_state145_133_1 + shifted_state145_133_3 + shifted_state145_133_5 + shifted_state145_145_0 + shifted_state145_145_1 + shifted_state145_145_2 + shifted_state145_145_5 + shifted_state145_145_6 + shifted_state145_145_7 + shifted_state145_153_1 + shifted_state145_167_0 + shifted_state145_167_1 + shifted_state145_167_2 + shifted_state145_167_5 + shifted_state145_181_0 + shifted_state145_181_2 + shifted_state145_181_3 + shifted_state145_181_4 + shifted_state145_181_5 + shifted_state145_181_6 + shifted_state145_181_7 + shifted_state145_186_3 + shifted_state145_186_4 + shifted_state145_187_0 + shifted_state145_187_1 + shifted_state145_187_2 + shifted_state145_187_5 + shifted_state145_187_6 + shifted_state145_187_7 + shifted_state145_188_1 + shifted_state145_188_3 + shifted_state145_188_4 + shifted_state145_188_6 + shifted_state145_188_7 + shifted_state145_189_3 + shifted_state145_189_4 + shifted_state145_199_1 + shifted_state145_199_2 + shifted_state145_199_3 + shifted_state145_199_4 + shifted_state145_199_5 + shifted_state145_199_6 + shifted_state145_199_7);
      reservoir_sum_parallel[146] = (shifted_state146_19_2 + shifted_state146_19_3 + shifted_state146_19_4 + shifted_state146_21_0 + shifted_state146_21_1 + shifted_state146_21_3 + shifted_state146_21_4 + shifted_state146_21_5 + shifted_state146_21_6 + shifted_state146_21_7 + shifted_state146_26_1 + shifted_state146_26_6 + shifted_state146_33_3 + shifted_state146_33_5 + shifted_state146_33_6 + shifted_state146_33_7 + shifted_state146_40_0 + shifted_state146_40_3 + shifted_state146_40_4 + shifted_state146_49_2 + shifted_state146_49_4 + shifted_state146_49_5 + shifted_state146_49_6 + shifted_state146_49_7 + shifted_state146_61_1 + shifted_state146_61_4 + shifted_state146_66_2 + shifted_state146_66_3 + shifted_state146_66_4 + shifted_state146_66_5 + shifted_state146_66_6 + shifted_state146_66_7 + shifted_state146_84_0 + shifted_state146_84_1 + shifted_state146_84_2 + shifted_state146_84_4 + shifted_state146_84_6 + shifted_state146_84_7 + shifted_state146_86_1 + shifted_state146_86_4 + shifted_state146_86_5 + shifted_state146_86_6 + shifted_state146_86_7 + shifted_state146_106_0 + shifted_state146_106_5 + shifted_state146_106_6 + shifted_state146_106_7 + shifted_state146_119_1 + shifted_state146_119_2 + shifted_state146_119_4 + shifted_state146_121_4 + shifted_state146_183_0 + shifted_state146_183_2 + shifted_state146_183_4 + shifted_state146_184_0 + shifted_state146_184_2 + shifted_state146_184_3 + shifted_state146_184_5 + shifted_state146_184_6 + shifted_state146_184_7 + shifted_state146_192_0 + shifted_state146_192_1 + shifted_state146_192_5 + shifted_state146_198_2);
      reservoir_sum_parallel[147] = (shifted_state147_21_0 + shifted_state147_21_1 + shifted_state147_21_4 + shifted_state147_29_3 + shifted_state147_29_4 + shifted_state147_50_1 + shifted_state147_50_2 + shifted_state147_50_3 + shifted_state147_50_5 + shifted_state147_50_6 + shifted_state147_50_7 + shifted_state147_59_1 + shifted_state147_59_2 + shifted_state147_59_3 + shifted_state147_59_4 + shifted_state147_59_5 + shifted_state147_59_6 + shifted_state147_59_7 + shifted_state147_60_0 + shifted_state147_60_1 + shifted_state147_60_2 + shifted_state147_60_3 + shifted_state147_60_5 + shifted_state147_60_6 + shifted_state147_60_7 + shifted_state147_66_0 + shifted_state147_66_1 + shifted_state147_66_4 + shifted_state147_66_5 + shifted_state147_66_6 + shifted_state147_66_7 + shifted_state147_93_1 + shifted_state147_93_2 + shifted_state147_93_3 + shifted_state147_93_5 + shifted_state147_93_6 + shifted_state147_93_7 + shifted_state147_95_2 + shifted_state147_95_3 + shifted_state147_97_1 + shifted_state147_97_2 + shifted_state147_97_3 + shifted_state147_97_4 + shifted_state147_135_0 + shifted_state147_135_1 + shifted_state147_135_2 + shifted_state147_135_3 + shifted_state147_135_5 + shifted_state147_141_0 + shifted_state147_141_1 + shifted_state147_141_2 + shifted_state147_147_0 + shifted_state147_147_1 + shifted_state147_147_4 + shifted_state147_147_5 + shifted_state147_147_6 + shifted_state147_147_7 + shifted_state147_160_1 + shifted_state147_160_3 + shifted_state147_160_5 + shifted_state147_160_6 + shifted_state147_160_7 + shifted_state147_178_0 + shifted_state147_178_3 + shifted_state147_178_5 + shifted_state147_178_6 + shifted_state147_178_7 + shifted_state147_183_2 + shifted_state147_183_3 + shifted_state147_183_5 + shifted_state147_183_6 + shifted_state147_183_7 + shifted_state147_190_1 + shifted_state147_190_4 + shifted_state147_190_5 + shifted_state147_190_6 + shifted_state147_190_7);
      reservoir_sum_parallel[148] = (shifted_state148_7_1 + shifted_state148_7_3 + shifted_state148_7_4 + shifted_state148_7_5 + shifted_state148_7_6 + shifted_state148_7_7 + shifted_state148_23_0 + shifted_state148_23_1 + shifted_state148_23_4 + shifted_state148_23_5 + shifted_state148_23_6 + shifted_state148_23_7 + shifted_state148_36_0 + shifted_state148_36_1 + shifted_state148_36_2 + shifted_state148_36_5 + shifted_state148_36_6 + shifted_state148_36_7 + shifted_state148_43_2 + shifted_state148_43_3 + shifted_state148_43_4 + shifted_state148_51_2 + shifted_state148_51_3 + shifted_state148_51_5 + shifted_state148_51_6 + shifted_state148_51_7 + shifted_state148_54_0 + shifted_state148_54_1 + shifted_state148_54_2 + shifted_state148_54_3 + shifted_state148_54_4 + shifted_state148_54_5 + shifted_state148_54_6 + shifted_state148_54_7 + shifted_state148_61_1 + shifted_state148_61_5 + shifted_state148_61_6 + shifted_state148_61_7 + shifted_state148_75_0 + shifted_state148_75_3 + shifted_state148_91_0 + shifted_state148_91_4 + shifted_state148_100_0 + shifted_state148_100_1 + shifted_state148_100_2 + shifted_state148_100_3 + shifted_state148_114_1 + shifted_state148_114_4 + shifted_state148_114_5 + shifted_state148_114_6 + shifted_state148_114_7 + shifted_state148_145_0 + shifted_state148_145_1 + shifted_state148_145_5 + shifted_state148_163_0 + shifted_state148_163_5 + shifted_state148_163_6 + shifted_state148_163_7 + shifted_state148_168_1 + shifted_state148_168_2 + shifted_state148_168_3 + shifted_state148_169_0 + shifted_state148_169_2 + shifted_state148_169_3 + shifted_state148_169_4 + shifted_state148_169_5 + shifted_state148_169_6 + shifted_state148_169_7 + shifted_state148_170_0 + shifted_state148_170_1 + shifted_state148_170_3 + shifted_state148_170_4 + shifted_state148_170_5 + shifted_state148_170_6 + shifted_state148_170_7 + shifted_state148_199_2 + shifted_state148_199_3 + shifted_state148_199_5 + shifted_state148_199_6 + shifted_state148_199_7);
      reservoir_sum_parallel[149] = (shifted_state149_6_4 + shifted_state149_6_5 + shifted_state149_6_6 + shifted_state149_6_7 + shifted_state149_62_3 + shifted_state149_63_1 + shifted_state149_63_2 + shifted_state149_63_3 + shifted_state149_63_5 + shifted_state149_63_6 + shifted_state149_63_7 + shifted_state149_83_1 + shifted_state149_83_3 + shifted_state149_100_1 + shifted_state149_100_3 + shifted_state149_100_6 + shifted_state149_100_7 + shifted_state149_103_4 + shifted_state149_123_1 + shifted_state149_123_2 + shifted_state149_123_5 + shifted_state149_136_0 + shifted_state149_136_1 + shifted_state149_136_4 + shifted_state149_136_5 + shifted_state149_136_6 + shifted_state149_136_7 + shifted_state149_149_2 + shifted_state149_149_3 + shifted_state149_149_4 + shifted_state149_149_6 + shifted_state149_149_7 + shifted_state149_159_0 + shifted_state149_159_4 + shifted_state149_159_5 + shifted_state149_160_0 + shifted_state149_160_1 + shifted_state149_160_2 + shifted_state149_160_4 + shifted_state149_166_1 + shifted_state149_166_4 + shifted_state149_166_5 + shifted_state149_166_6 + shifted_state149_166_7 + shifted_state149_167_1 + shifted_state149_167_3 + shifted_state149_167_4 + shifted_state149_172_0 + shifted_state149_172_1 + shifted_state149_172_4 + shifted_state149_172_6 + shifted_state149_172_7 + shifted_state149_174_1 + shifted_state149_174_2 + shifted_state149_174_3 + shifted_state149_174_5 + shifted_state149_174_7);
      reservoir_sum_parallel[150] = (shifted_state150_7_0 + shifted_state150_7_1 + shifted_state150_7_2 + shifted_state150_7_5 + shifted_state150_7_6 + shifted_state150_7_7 + shifted_state150_12_2 + shifted_state150_12_3 + shifted_state150_12_5 + shifted_state150_12_6 + shifted_state150_12_7 + shifted_state150_21_1 + shifted_state150_21_2 + shifted_state150_21_3 + shifted_state150_21_4 + shifted_state150_21_5 + shifted_state150_21_6 + shifted_state150_21_7 + shifted_state150_41_0 + shifted_state150_41_1 + shifted_state150_41_2 + shifted_state150_45_0 + shifted_state150_45_3 + shifted_state150_45_4 + shifted_state150_45_5 + shifted_state150_45_6 + shifted_state150_45_7 + shifted_state150_54_3 + shifted_state150_54_4 + shifted_state150_54_5 + shifted_state150_54_6 + shifted_state150_54_7 + shifted_state150_59_0 + shifted_state150_59_1 + shifted_state150_60_0 + shifted_state150_60_1 + shifted_state150_60_2 + shifted_state150_60_3 + shifted_state150_60_4 + shifted_state150_60_5 + shifted_state150_62_0 + shifted_state150_62_5 + shifted_state150_62_6 + shifted_state150_62_7 + shifted_state150_68_0 + shifted_state150_68_2 + shifted_state150_68_5 + shifted_state150_94_4 + shifted_state150_94_5 + shifted_state150_94_6 + shifted_state150_94_7 + shifted_state150_109_1 + shifted_state150_109_6 + shifted_state150_109_7 + shifted_state150_113_0 + shifted_state150_113_2 + shifted_state150_129_1 + shifted_state150_129_2 + shifted_state150_129_5 + shifted_state150_129_6 + shifted_state150_129_7 + shifted_state150_132_0 + shifted_state150_132_3 + shifted_state150_132_4 + shifted_state150_132_5 + shifted_state150_132_6 + shifted_state150_132_7 + shifted_state150_136_0 + shifted_state150_136_3 + shifted_state150_141_1 + shifted_state150_141_2 + shifted_state150_141_5 + shifted_state150_148_1 + shifted_state150_148_4 + shifted_state150_161_1 + shifted_state150_161_3 + shifted_state150_161_4 + shifted_state150_162_3 + shifted_state150_162_5 + shifted_state150_163_6 + shifted_state150_163_7 + shifted_state150_164_0 + shifted_state150_164_1 + shifted_state150_164_2 + shifted_state150_164_4 + shifted_state150_170_1 + shifted_state150_170_5 + shifted_state150_170_6 + shifted_state150_170_7 + shifted_state150_178_0 + shifted_state150_178_1 + shifted_state150_178_2 + shifted_state150_178_3 + shifted_state150_199_1 + shifted_state150_199_5 + shifted_state150_199_6 + shifted_state150_199_7);
      reservoir_sum_parallel[151] = (shifted_state151_6_0 + shifted_state151_6_3 + shifted_state151_7_0 + shifted_state151_7_1 + shifted_state151_7_5 + shifted_state151_7_6 + shifted_state151_7_7 + shifted_state151_18_1 + shifted_state151_18_2 + shifted_state151_18_3 + shifted_state151_32_3 + shifted_state151_32_4 + shifted_state151_43_2 + shifted_state151_43_4 + shifted_state151_62_1 + shifted_state151_62_2 + shifted_state151_62_4 + shifted_state151_62_5 + shifted_state151_62_6 + shifted_state151_62_7 + shifted_state151_92_2 + shifted_state151_92_3 + shifted_state151_92_4 + shifted_state151_92_5 + shifted_state151_92_6 + shifted_state151_92_7 + shifted_state151_94_0 + shifted_state151_94_3 + shifted_state151_94_6 + shifted_state151_94_7 + shifted_state151_115_0 + shifted_state151_115_1 + shifted_state151_115_5 + shifted_state151_115_6 + shifted_state151_115_7 + shifted_state151_116_0 + shifted_state151_116_1 + shifted_state151_116_3 + shifted_state151_116_5 + shifted_state151_116_6 + shifted_state151_116_7 + shifted_state151_124_0 + shifted_state151_124_1 + shifted_state151_124_2 + shifted_state151_124_3 + shifted_state151_124_4 + shifted_state151_124_5 + shifted_state151_124_6 + shifted_state151_124_7 + shifted_state151_130_0 + shifted_state151_130_1 + shifted_state151_130_2 + shifted_state151_130_3 + shifted_state151_130_5 + shifted_state151_130_6 + shifted_state151_130_7 + shifted_state151_133_1 + shifted_state151_133_2 + shifted_state151_133_3 + shifted_state151_133_4 + shifted_state151_133_5 + shifted_state151_133_6 + shifted_state151_133_7 + shifted_state151_157_1 + shifted_state151_157_4 + shifted_state151_157_5 + shifted_state151_178_0 + shifted_state151_178_2 + shifted_state151_178_3 + shifted_state151_178_4 + shifted_state151_178_6 + shifted_state151_178_7 + shifted_state151_180_0 + shifted_state151_180_1 + shifted_state151_180_2);
      reservoir_sum_parallel[152] = (shifted_state152_5_1 + shifted_state152_5_2 + shifted_state152_5_6 + shifted_state152_5_7 + shifted_state152_11_0 + shifted_state152_11_1 + shifted_state152_11_3 + shifted_state152_11_5 + shifted_state152_11_6 + shifted_state152_11_7 + shifted_state152_22_0 + shifted_state152_22_1 + shifted_state152_22_4 + shifted_state152_35_0 + shifted_state152_35_2 + shifted_state152_35_4 + shifted_state152_35_6 + shifted_state152_35_7 + shifted_state152_47_0 + shifted_state152_47_2 + shifted_state152_47_3 + shifted_state152_47_4 + shifted_state152_47_6 + shifted_state152_47_7 + shifted_state152_52_0 + shifted_state152_52_3 + shifted_state152_66_0 + shifted_state152_66_2 + shifted_state152_66_6 + shifted_state152_72_1 + shifted_state152_72_2 + shifted_state152_72_3 + shifted_state152_72_4 + shifted_state152_72_5 + shifted_state152_72_6 + shifted_state152_72_7 + shifted_state152_86_0 + shifted_state152_86_1 + shifted_state152_86_3 + shifted_state152_86_4 + shifted_state152_86_5 + shifted_state152_86_6 + shifted_state152_86_7 + shifted_state152_90_0 + shifted_state152_100_0 + shifted_state152_100_1 + shifted_state152_100_3 + shifted_state152_100_4 + shifted_state152_100_5 + shifted_state152_100_7 + shifted_state152_101_5 + shifted_state152_101_6 + shifted_state152_101_7 + shifted_state152_102_1 + shifted_state152_102_3 + shifted_state152_102_6 + shifted_state152_116_0 + shifted_state152_116_2 + shifted_state152_116_3 + shifted_state152_116_4 + shifted_state152_116_6 + shifted_state152_116_7 + shifted_state152_139_0 + shifted_state152_139_2 + shifted_state152_139_4 + shifted_state152_139_5 + shifted_state152_139_6 + shifted_state152_139_7 + shifted_state152_152_1 + shifted_state152_152_2 + shifted_state152_152_4 + shifted_state152_159_3 + shifted_state152_195_0 + shifted_state152_195_2);
      reservoir_sum_parallel[153] = (shifted_state153_15_1 + shifted_state153_15_5 + shifted_state153_15_6 + shifted_state153_15_7 + shifted_state153_18_0 + shifted_state153_18_2 + shifted_state153_18_4 + shifted_state153_18_6 + shifted_state153_18_7 + shifted_state153_22_1 + shifted_state153_22_3 + shifted_state153_22_4 + shifted_state153_22_6 + shifted_state153_22_7 + shifted_state153_28_2 + shifted_state153_28_4 + shifted_state153_28_5 + shifted_state153_28_6 + shifted_state153_28_7 + shifted_state153_44_1 + shifted_state153_44_3 + shifted_state153_44_5 + shifted_state153_44_6 + shifted_state153_44_7 + shifted_state153_46_3 + shifted_state153_46_4 + shifted_state153_46_5 + shifted_state153_46_6 + shifted_state153_46_7 + shifted_state153_62_0 + shifted_state153_62_2 + shifted_state153_62_3 + shifted_state153_62_4 + shifted_state153_73_3 + shifted_state153_73_4 + shifted_state153_73_5 + shifted_state153_73_6 + shifted_state153_73_7 + shifted_state153_75_0 + shifted_state153_75_4 + shifted_state153_75_5 + shifted_state153_75_6 + shifted_state153_75_7 + shifted_state153_91_3 + shifted_state153_91_5 + shifted_state153_91_6 + shifted_state153_91_7 + shifted_state153_93_0 + shifted_state153_93_1 + shifted_state153_93_2 + shifted_state153_93_3 + shifted_state153_93_6 + shifted_state153_93_7 + shifted_state153_104_2 + shifted_state153_104_3 + shifted_state153_104_5 + shifted_state153_104_6 + shifted_state153_104_7 + shifted_state153_108_2 + shifted_state153_108_3 + shifted_state153_108_4 + shifted_state153_108_5 + shifted_state153_108_6 + shifted_state153_108_7 + shifted_state153_113_1 + shifted_state153_113_2 + shifted_state153_113_3 + shifted_state153_113_4 + shifted_state153_113_5 + shifted_state153_113_6 + shifted_state153_113_7 + shifted_state153_118_2 + shifted_state153_122_2 + shifted_state153_129_0 + shifted_state153_129_2 + shifted_state153_129_3 + shifted_state153_129_4 + shifted_state153_129_6 + shifted_state153_129_7 + shifted_state153_130_3 + shifted_state153_130_4 + shifted_state153_130_5 + shifted_state153_140_2 + shifted_state153_140_3 + shifted_state153_140_4 + shifted_state153_140_5 + shifted_state153_140_6 + shifted_state153_140_7 + shifted_state153_150_0 + shifted_state153_150_1 + shifted_state153_150_2 + shifted_state153_150_3 + shifted_state153_150_4 + shifted_state153_150_5 + shifted_state153_150_7 + shifted_state153_152_1 + shifted_state153_152_4 + shifted_state153_152_5 + shifted_state153_152_6 + shifted_state153_152_7 + shifted_state153_164_4 + shifted_state153_164_6 + shifted_state153_164_7 + shifted_state153_165_0 + shifted_state153_165_2 + shifted_state153_165_3 + shifted_state153_165_4 + shifted_state153_165_5 + shifted_state153_165_6 + shifted_state153_165_7 + shifted_state153_184_1 + shifted_state153_184_2 + shifted_state153_184_3 + shifted_state153_184_5 + shifted_state153_184_6 + shifted_state153_184_7);
      reservoir_sum_parallel[154] = (shifted_state154_8_0 + shifted_state154_8_1 + shifted_state154_8_2 + shifted_state154_8_3 + shifted_state154_31_3 + shifted_state154_31_6 + shifted_state154_31_7 + shifted_state154_37_1 + shifted_state154_37_2 + shifted_state154_37_3 + shifted_state154_37_5 + shifted_state154_37_6 + shifted_state154_37_7 + shifted_state154_50_2 + shifted_state154_50_3 + shifted_state154_50_6 + shifted_state154_50_7 + shifted_state154_53_2 + shifted_state154_53_3 + shifted_state154_53_5 + shifted_state154_53_6 + shifted_state154_53_7 + shifted_state154_59_1 + shifted_state154_59_2 + shifted_state154_59_3 + shifted_state154_59_5 + shifted_state154_59_6 + shifted_state154_59_7 + shifted_state154_69_0 + shifted_state154_69_3 + shifted_state154_69_4 + shifted_state154_78_0 + shifted_state154_78_1 + shifted_state154_78_3 + shifted_state154_78_5 + shifted_state154_85_2 + shifted_state154_89_0 + shifted_state154_89_3 + shifted_state154_89_4 + shifted_state154_89_5 + shifted_state154_89_6 + shifted_state154_89_7 + shifted_state154_99_2 + shifted_state154_99_4 + shifted_state154_99_5 + shifted_state154_99_6 + shifted_state154_99_7 + shifted_state154_114_0 + shifted_state154_114_3 + shifted_state154_114_4 + shifted_state154_114_5 + shifted_state154_114_6 + shifted_state154_114_7 + shifted_state154_125_0 + shifted_state154_125_1 + shifted_state154_125_2 + shifted_state154_125_3 + shifted_state154_125_5 + shifted_state154_125_6 + shifted_state154_125_7 + shifted_state154_157_2 + shifted_state154_157_3 + shifted_state154_171_5 + shifted_state154_171_6 + shifted_state154_171_7 + shifted_state154_172_1 + shifted_state154_172_2 + shifted_state154_172_3 + shifted_state154_172_4 + shifted_state154_172_5 + shifted_state154_172_6 + shifted_state154_172_7 + shifted_state154_177_2 + shifted_state154_177_3 + shifted_state154_177_4 + shifted_state154_187_0 + shifted_state154_187_3 + shifted_state154_187_4);
      reservoir_sum_parallel[155] = (shifted_state155_4_1 + shifted_state155_4_2 + shifted_state155_4_3 + shifted_state155_4_5 + shifted_state155_4_6 + shifted_state155_4_7 + shifted_state155_7_0 + shifted_state155_7_1 + shifted_state155_7_4 + shifted_state155_7_5 + shifted_state155_7_6 + shifted_state155_7_7 + shifted_state155_11_1 + shifted_state155_11_4 + shifted_state155_16_0 + shifted_state155_16_1 + shifted_state155_16_3 + shifted_state155_16_4 + shifted_state155_17_0 + shifted_state155_17_1 + shifted_state155_17_5 + shifted_state155_17_6 + shifted_state155_17_7 + shifted_state155_60_1 + shifted_state155_60_3 + shifted_state155_61_0 + shifted_state155_61_1 + shifted_state155_61_3 + shifted_state155_61_4 + shifted_state155_61_5 + shifted_state155_61_6 + shifted_state155_61_7 + shifted_state155_71_3 + shifted_state155_72_0 + shifted_state155_72_1 + shifted_state155_72_3 + shifted_state155_92_0 + shifted_state155_92_1 + shifted_state155_92_3 + shifted_state155_97_0 + shifted_state155_97_3 + shifted_state155_97_4 + shifted_state155_97_5 + shifted_state155_97_6 + shifted_state155_97_7 + shifted_state155_107_2 + shifted_state155_107_3 + shifted_state155_107_5 + shifted_state155_107_6 + shifted_state155_107_7 + shifted_state155_125_1 + shifted_state155_125_5 + shifted_state155_125_6 + shifted_state155_125_7 + shifted_state155_131_0 + shifted_state155_131_4 + shifted_state155_142_1 + shifted_state155_142_2 + shifted_state155_142_3 + shifted_state155_148_0 + shifted_state155_148_2 + shifted_state155_149_0 + shifted_state155_149_4 + shifted_state155_155_0 + shifted_state155_155_2 + shifted_state155_155_3 + shifted_state155_155_5 + shifted_state155_155_6 + shifted_state155_155_7 + shifted_state155_164_0 + shifted_state155_164_3 + shifted_state155_164_4 + shifted_state155_164_5 + shifted_state155_164_6 + shifted_state155_164_7 + shifted_state155_168_2 + shifted_state155_168_4 + shifted_state155_186_1 + shifted_state155_186_3 + shifted_state155_186_5 + shifted_state155_186_6 + shifted_state155_186_7 + shifted_state155_190_0 + shifted_state155_190_3 + shifted_state155_190_5 + shifted_state155_190_6 + shifted_state155_190_7 + shifted_state155_193_2 + shifted_state155_193_3 + shifted_state155_193_5 + shifted_state155_193_6 + shifted_state155_193_7 + shifted_state155_194_0 + shifted_state155_194_1 + shifted_state155_194_2 + shifted_state155_194_3 + shifted_state155_194_4 + shifted_state155_194_5);
      reservoir_sum_parallel[156] = (shifted_state156_4_1 + shifted_state156_4_2 + shifted_state156_4_4 + shifted_state156_5_1 + shifted_state156_5_2 + shifted_state156_17_0 + shifted_state156_17_1 + shifted_state156_17_3 + shifted_state156_20_0 + shifted_state156_20_1 + shifted_state156_20_2 + shifted_state156_20_3 + shifted_state156_20_4 + shifted_state156_20_5 + shifted_state156_20_6 + shifted_state156_20_7 + shifted_state156_31_0 + shifted_state156_31_1 + shifted_state156_31_3 + shifted_state156_35_1 + shifted_state156_38_0 + shifted_state156_38_2 + shifted_state156_38_3 + shifted_state156_38_5 + shifted_state156_38_6 + shifted_state156_38_7 + shifted_state156_40_1 + shifted_state156_40_2 + shifted_state156_40_3 + shifted_state156_40_4 + shifted_state156_40_6 + shifted_state156_40_7 + shifted_state156_43_0 + shifted_state156_43_1 + shifted_state156_43_2 + shifted_state156_43_3 + shifted_state156_44_0 + shifted_state156_44_1 + shifted_state156_44_2 + shifted_state156_44_3 + shifted_state156_44_4 + shifted_state156_44_5 + shifted_state156_44_6 + shifted_state156_44_7 + shifted_state156_47_0 + shifted_state156_47_3 + shifted_state156_55_4 + shifted_state156_63_0 + shifted_state156_63_2 + shifted_state156_63_3 + shifted_state156_80_1 + shifted_state156_80_2 + shifted_state156_80_3 + shifted_state156_80_4 + shifted_state156_107_0 + shifted_state156_107_1 + shifted_state156_107_3 + shifted_state156_150_0 + shifted_state156_150_3 + shifted_state156_150_4 + shifted_state156_150_5 + shifted_state156_150_6 + shifted_state156_150_7 + shifted_state156_168_0 + shifted_state156_168_1 + shifted_state156_168_3 + shifted_state156_168_4 + shifted_state156_168_6 + shifted_state156_168_7 + shifted_state156_177_2 + shifted_state156_177_3 + shifted_state156_177_4 + shifted_state156_177_5 + shifted_state156_177_6 + shifted_state156_177_7 + shifted_state156_183_0 + shifted_state156_183_3 + shifted_state156_183_5 + shifted_state156_183_6 + shifted_state156_183_7 + shifted_state156_192_0 + shifted_state156_192_4 + shifted_state156_194_0 + shifted_state156_194_1 + shifted_state156_194_2 + shifted_state156_194_3 + shifted_state156_194_4 + shifted_state156_194_5 + shifted_state156_194_6 + shifted_state156_194_7 + shifted_state156_198_0 + shifted_state156_198_1 + shifted_state156_198_3 + shifted_state156_198_4 + shifted_state156_198_5 + shifted_state156_198_6 + shifted_state156_198_7);
      reservoir_sum_parallel[157] = (shifted_state157_9_1 + shifted_state157_9_5 + shifted_state157_10_3 + shifted_state157_10_5 + shifted_state157_10_6 + shifted_state157_10_7 + shifted_state157_24_1 + shifted_state157_24_3 + shifted_state157_24_5 + shifted_state157_30_1 + shifted_state157_30_4 + shifted_state157_31_0 + shifted_state157_31_4 + shifted_state157_32_3 + shifted_state157_32_4 + shifted_state157_32_5 + shifted_state157_32_6 + shifted_state157_32_7 + shifted_state157_50_1 + shifted_state157_50_2 + shifted_state157_50_3 + shifted_state157_50_5 + shifted_state157_50_6 + shifted_state157_50_7 + shifted_state157_86_1 + shifted_state157_86_3 + shifted_state157_86_5 + shifted_state157_86_6 + shifted_state157_86_7 + shifted_state157_87_1 + shifted_state157_87_4 + shifted_state157_87_5 + shifted_state157_87_6 + shifted_state157_87_7 + shifted_state157_96_2 + shifted_state157_103_1 + shifted_state157_103_2 + shifted_state157_103_3 + shifted_state157_113_1 + shifted_state157_113_2 + shifted_state157_113_4 + shifted_state157_117_3 + shifted_state157_117_5 + shifted_state157_117_6 + shifted_state157_117_7 + shifted_state157_123_0 + shifted_state157_123_5 + shifted_state157_133_0 + shifted_state157_133_1 + shifted_state157_133_4 + shifted_state157_135_0 + shifted_state157_135_2 + shifted_state157_154_0 + shifted_state157_154_3 + shifted_state157_154_4 + shifted_state157_154_5 + shifted_state157_154_6 + shifted_state157_154_7 + shifted_state157_155_0 + shifted_state157_155_3);
      reservoir_sum_parallel[158] = (shifted_state158_3_2 + shifted_state158_3_3 + shifted_state158_3_4 + shifted_state158_3_5 + shifted_state158_3_6 + shifted_state158_3_7 + shifted_state158_15_2 + shifted_state158_15_5 + shifted_state158_25_2 + shifted_state158_25_3 + shifted_state158_25_4 + shifted_state158_25_5 + shifted_state158_25_6 + shifted_state158_25_7 + shifted_state158_50_3 + shifted_state158_50_5 + shifted_state158_50_6 + shifted_state158_50_7 + shifted_state158_58_0 + shifted_state158_58_1 + shifted_state158_58_3 + shifted_state158_58_5 + shifted_state158_58_6 + shifted_state158_58_7 + shifted_state158_60_1 + shifted_state158_60_5 + shifted_state158_60_6 + shifted_state158_60_7 + shifted_state158_67_1 + shifted_state158_82_0 + shifted_state158_82_1 + shifted_state158_82_2 + shifted_state158_86_0 + shifted_state158_86_1 + shifted_state158_86_2 + shifted_state158_86_3 + shifted_state158_86_4 + shifted_state158_86_5 + shifted_state158_86_6 + shifted_state158_86_7 + shifted_state158_89_0 + shifted_state158_89_2 + shifted_state158_89_4 + shifted_state158_89_5 + shifted_state158_89_6 + shifted_state158_89_7 + shifted_state158_113_0 + shifted_state158_113_2 + shifted_state158_113_3 + shifted_state158_114_0 + shifted_state158_114_1 + shifted_state158_145_0 + shifted_state158_145_1 + shifted_state158_145_2 + shifted_state158_145_4 + shifted_state158_160_3 + shifted_state158_160_4 + shifted_state158_160_6 + shifted_state158_160_7 + shifted_state158_171_0 + shifted_state158_171_1 + shifted_state158_171_2 + shifted_state158_171_4 + shifted_state158_177_4 + shifted_state158_185_4 + shifted_state158_185_5 + shifted_state158_185_6 + shifted_state158_185_7 + shifted_state158_190_0 + shifted_state158_190_2 + shifted_state158_190_3 + shifted_state158_190_4 + shifted_state158_195_0 + shifted_state158_195_3 + shifted_state158_195_5);
      reservoir_sum_parallel[159] = (shifted_state159_0_2 + shifted_state159_0_3 + shifted_state159_0_5 + shifted_state159_0_6 + shifted_state159_0_7 + shifted_state159_14_1 + shifted_state159_14_4 + shifted_state159_14_5 + shifted_state159_14_6 + shifted_state159_14_7 + shifted_state159_21_1 + shifted_state159_21_2 + shifted_state159_37_0 + shifted_state159_37_3 + shifted_state159_37_4 + shifted_state159_48_0 + shifted_state159_48_1 + shifted_state159_48_2 + shifted_state159_51_1 + shifted_state159_51_6 + shifted_state159_64_0 + shifted_state159_64_3 + shifted_state159_105_0 + shifted_state159_116_0 + shifted_state159_116_1 + shifted_state159_116_2 + shifted_state159_116_3 + shifted_state159_116_4 + shifted_state159_116_6 + shifted_state159_116_7 + shifted_state159_140_1 + shifted_state159_140_2 + shifted_state159_140_5 + shifted_state159_141_1 + shifted_state159_141_4 + shifted_state159_146_1 + shifted_state159_146_2 + shifted_state159_146_3 + shifted_state159_146_4 + shifted_state159_146_6 + shifted_state159_146_7 + shifted_state159_154_0 + shifted_state159_154_2 + shifted_state159_154_4 + shifted_state159_154_5 + shifted_state159_154_6 + shifted_state159_154_7 + shifted_state159_182_0 + shifted_state159_182_2 + shifted_state159_182_3 + shifted_state159_182_4 + shifted_state159_182_5 + shifted_state159_182_6 + shifted_state159_182_7);
      reservoir_sum_parallel[160] = (shifted_state160_16_1 + shifted_state160_16_2 + shifted_state160_16_5 + shifted_state160_16_6 + shifted_state160_16_7 + shifted_state160_29_0 + shifted_state160_29_4 + shifted_state160_29_6 + shifted_state160_29_7 + shifted_state160_33_2 + shifted_state160_33_4 + shifted_state160_47_1 + shifted_state160_47_3 + shifted_state160_47_4 + shifted_state160_47_6 + shifted_state160_47_7 + shifted_state160_55_1 + shifted_state160_55_3 + shifted_state160_55_5 + shifted_state160_56_3 + shifted_state160_56_4 + shifted_state160_56_5 + shifted_state160_56_6 + shifted_state160_56_7 + shifted_state160_59_1 + shifted_state160_59_2 + shifted_state160_59_3 + shifted_state160_69_0 + shifted_state160_69_2 + shifted_state160_69_3 + shifted_state160_69_4 + shifted_state160_72_3 + shifted_state160_72_5 + shifted_state160_72_6 + shifted_state160_72_7 + shifted_state160_79_4 + shifted_state160_82_1 + shifted_state160_82_2 + shifted_state160_82_4 + shifted_state160_82_6 + shifted_state160_82_7 + shifted_state160_103_1 + shifted_state160_103_3 + shifted_state160_103_4 + shifted_state160_104_0 + shifted_state160_104_1 + shifted_state160_104_2 + shifted_state160_104_3 + shifted_state160_105_1 + shifted_state160_105_2 + shifted_state160_105_4 + shifted_state160_105_5 + shifted_state160_105_6 + shifted_state160_105_7 + shifted_state160_113_0 + shifted_state160_113_1 + shifted_state160_113_4 + shifted_state160_117_1 + shifted_state160_117_2 + shifted_state160_117_3 + shifted_state160_118_2 + shifted_state160_118_3 + shifted_state160_119_4 + shifted_state160_124_3 + shifted_state160_157_1 + shifted_state160_157_2 + shifted_state160_157_4 + shifted_state160_157_5 + shifted_state160_157_6 + shifted_state160_157_7 + shifted_state160_158_2 + shifted_state160_158_4 + shifted_state160_163_0 + shifted_state160_163_5 + shifted_state160_170_3 + shifted_state160_170_4 + shifted_state160_170_5 + shifted_state160_170_6 + shifted_state160_170_7);
      reservoir_sum_parallel[161] = (shifted_state161_27_0 + shifted_state161_27_1 + shifted_state161_43_0 + shifted_state161_43_3 + shifted_state161_43_4 + shifted_state161_43_6 + shifted_state161_43_7 + shifted_state161_48_0 + shifted_state161_48_1 + shifted_state161_48_2 + shifted_state161_48_3 + shifted_state161_48_4 + shifted_state161_65_0 + shifted_state161_65_1 + shifted_state161_65_3 + shifted_state161_65_4 + shifted_state161_65_5 + shifted_state161_65_6 + shifted_state161_65_7 + shifted_state161_73_4 + shifted_state161_76_4 + shifted_state161_85_1 + shifted_state161_85_2 + shifted_state161_85_4 + shifted_state161_85_5 + shifted_state161_85_6 + shifted_state161_85_7 + shifted_state161_87_0 + shifted_state161_87_4 + shifted_state161_87_5 + shifted_state161_87_6 + shifted_state161_87_7 + shifted_state161_111_1 + shifted_state161_111_2 + shifted_state161_111_4 + shifted_state161_111_5 + shifted_state161_111_6 + shifted_state161_111_7 + shifted_state161_113_0 + shifted_state161_113_2 + shifted_state161_113_4 + shifted_state161_113_5 + shifted_state161_113_6 + shifted_state161_113_7 + shifted_state161_124_0 + shifted_state161_124_1 + shifted_state161_124_4 + shifted_state161_124_5 + shifted_state161_124_7 + shifted_state161_137_1 + shifted_state161_137_3 + shifted_state161_137_5 + shifted_state161_137_6 + shifted_state161_137_7 + shifted_state161_152_1 + shifted_state161_152_2 + shifted_state161_152_5 + shifted_state161_152_6 + shifted_state161_152_7 + shifted_state161_161_0 + shifted_state161_161_2 + shifted_state161_161_4 + shifted_state161_161_6 + shifted_state161_161_7 + shifted_state161_187_3 + shifted_state161_187_6);
      reservoir_sum_parallel[162] = (shifted_state162_9_3 + shifted_state162_9_4 + shifted_state162_13_1 + shifted_state162_13_2 + shifted_state162_13_4 + shifted_state162_13_6 + shifted_state162_13_7 + shifted_state162_21_1 + shifted_state162_21_3 + shifted_state162_21_4 + shifted_state162_21_5 + shifted_state162_21_6 + shifted_state162_21_7 + shifted_state162_25_0 + shifted_state162_25_1 + shifted_state162_25_2 + shifted_state162_25_3 + shifted_state162_25_4 + shifted_state162_26_3 + shifted_state162_26_5 + shifted_state162_31_3 + shifted_state162_31_4 + shifted_state162_31_5 + shifted_state162_31_6 + shifted_state162_31_7 + shifted_state162_40_0 + shifted_state162_40_2 + shifted_state162_40_3 + shifted_state162_40_4 + shifted_state162_40_5 + shifted_state162_40_6 + shifted_state162_40_7 + shifted_state162_55_2 + shifted_state162_55_4 + shifted_state162_55_5 + shifted_state162_55_6 + shifted_state162_55_7 + shifted_state162_58_0 + shifted_state162_58_3 + shifted_state162_58_4 + shifted_state162_59_0 + shifted_state162_59_1 + shifted_state162_92_0 + shifted_state162_92_4 + shifted_state162_92_5 + shifted_state162_96_1 + shifted_state162_96_3 + shifted_state162_96_4 + shifted_state162_96_5 + shifted_state162_96_6 + shifted_state162_96_7 + shifted_state162_102_0 + shifted_state162_102_4 + shifted_state162_102_5 + shifted_state162_102_6 + shifted_state162_102_7 + shifted_state162_132_0 + shifted_state162_132_1 + shifted_state162_132_3 + shifted_state162_132_4 + shifted_state162_132_6 + shifted_state162_132_7 + shifted_state162_143_4 + shifted_state162_143_5 + shifted_state162_143_6 + shifted_state162_143_7 + shifted_state162_149_0 + shifted_state162_149_1 + shifted_state162_149_4 + shifted_state162_149_5 + shifted_state162_149_6 + shifted_state162_149_7 + shifted_state162_155_0 + shifted_state162_155_3);
      reservoir_sum_parallel[163] = (shifted_state163_4_1 + shifted_state163_4_3 + shifted_state163_24_4 + shifted_state163_45_2 + shifted_state163_45_5 + shifted_state163_45_6 + shifted_state163_45_7 + shifted_state163_52_0 + shifted_state163_52_1 + shifted_state163_63_0 + shifted_state163_63_1 + shifted_state163_63_2 + shifted_state163_71_0 + shifted_state163_71_3 + shifted_state163_71_4 + shifted_state163_71_6 + shifted_state163_71_7 + shifted_state163_78_1 + shifted_state163_78_3 + shifted_state163_78_4 + shifted_state163_78_6 + shifted_state163_78_7 + shifted_state163_81_3 + shifted_state163_81_5 + shifted_state163_81_6 + shifted_state163_81_7 + shifted_state163_94_0 + shifted_state163_94_1 + shifted_state163_94_5 + shifted_state163_94_6 + shifted_state163_94_7 + shifted_state163_98_0 + shifted_state163_98_1 + shifted_state163_98_2 + shifted_state163_98_3 + shifted_state163_98_4 + shifted_state163_145_2 + shifted_state163_145_5 + shifted_state163_145_6 + shifted_state163_145_7 + shifted_state163_175_1 + shifted_state163_175_6 + shifted_state163_175_7 + shifted_state163_178_0 + shifted_state163_178_2 + shifted_state163_178_4 + shifted_state163_178_5 + shifted_state163_178_6 + shifted_state163_178_7 + shifted_state163_182_0 + shifted_state163_182_4 + shifted_state163_182_5 + shifted_state163_182_6 + shifted_state163_182_7 + shifted_state163_187_0 + shifted_state163_187_1 + shifted_state163_187_2 + shifted_state163_187_4 + shifted_state163_192_0 + shifted_state163_192_1 + shifted_state163_192_3 + shifted_state163_192_5 + shifted_state163_192_6 + shifted_state163_192_7 + shifted_state163_193_1 + shifted_state163_193_2 + shifted_state163_193_3 + shifted_state163_194_0 + shifted_state163_194_3 + shifted_state163_194_6 + shifted_state163_194_7 + shifted_state163_196_4 + shifted_state163_196_5 + shifted_state163_196_6 + shifted_state163_196_7 + shifted_state163_197_0 + shifted_state163_197_1 + shifted_state163_197_4);
      reservoir_sum_parallel[164] = (shifted_state164_2_1 + shifted_state164_2_4 + shifted_state164_10_0 + shifted_state164_10_3 + shifted_state164_10_6 + shifted_state164_11_0 + shifted_state164_11_2 + shifted_state164_11_3 + shifted_state164_11_5 + shifted_state164_13_0 + shifted_state164_13_2 + shifted_state164_13_4 + shifted_state164_13_5 + shifted_state164_13_6 + shifted_state164_13_7 + shifted_state164_18_0 + shifted_state164_18_2 + shifted_state164_18_5 + shifted_state164_18_6 + shifted_state164_18_7 + shifted_state164_20_2 + shifted_state164_20_3 + shifted_state164_20_4 + shifted_state164_29_0 + shifted_state164_29_4 + shifted_state164_29_5 + shifted_state164_32_0 + shifted_state164_32_1 + shifted_state164_32_4 + shifted_state164_32_5 + shifted_state164_39_1 + shifted_state164_39_2 + shifted_state164_39_3 + shifted_state164_39_4 + shifted_state164_39_5 + shifted_state164_39_6 + shifted_state164_39_7 + shifted_state164_47_0 + shifted_state164_47_1 + shifted_state164_47_2 + shifted_state164_47_4 + shifted_state164_47_5 + shifted_state164_47_6 + shifted_state164_47_7 + shifted_state164_54_1 + shifted_state164_54_2 + shifted_state164_54_3 + shifted_state164_54_5 + shifted_state164_54_6 + shifted_state164_54_7 + shifted_state164_69_0 + shifted_state164_69_2 + shifted_state164_69_4 + shifted_state164_69_5 + shifted_state164_69_6 + shifted_state164_69_7 + shifted_state164_77_1 + shifted_state164_77_2 + shifted_state164_77_3 + shifted_state164_77_4 + shifted_state164_77_5 + shifted_state164_77_6 + shifted_state164_77_7 + shifted_state164_85_0 + shifted_state164_85_1 + shifted_state164_85_2 + shifted_state164_88_1 + shifted_state164_88_3 + shifted_state164_88_4 + shifted_state164_89_1 + shifted_state164_89_3 + shifted_state164_89_4 + shifted_state164_89_6 + shifted_state164_94_0 + shifted_state164_94_1 + shifted_state164_94_3 + shifted_state164_94_5 + shifted_state164_115_1 + shifted_state164_115_2 + shifted_state164_116_0 + shifted_state164_116_3 + shifted_state164_116_4 + shifted_state164_122_0 + shifted_state164_122_2 + shifted_state164_122_3 + shifted_state164_122_4 + shifted_state164_122_6 + shifted_state164_122_7 + shifted_state164_130_1 + shifted_state164_130_2 + shifted_state164_130_3 + shifted_state164_130_4 + shifted_state164_133_0 + shifted_state164_133_2 + shifted_state164_133_4 + shifted_state164_140_3 + shifted_state164_154_0 + shifted_state164_154_1 + shifted_state164_154_2 + shifted_state164_154_3 + shifted_state164_154_5 + shifted_state164_188_2 + shifted_state164_188_4 + shifted_state164_188_5 + shifted_state164_192_1 + shifted_state164_192_2 + shifted_state164_192_3 + shifted_state164_192_4 + shifted_state164_192_5 + shifted_state164_192_6 + shifted_state164_192_7 + shifted_state164_193_4 + shifted_state164_193_5 + shifted_state164_193_6 + shifted_state164_193_7 + shifted_state164_194_3 + shifted_state164_194_5 + shifted_state164_194_6 + shifted_state164_194_7);
      reservoir_sum_parallel[165] = (shifted_state165_13_1 + shifted_state165_13_2 + shifted_state165_13_3 + shifted_state165_13_5 + shifted_state165_13_6 + shifted_state165_13_7 + shifted_state165_27_0 + shifted_state165_27_3 + shifted_state165_27_4 + shifted_state165_74_2 + shifted_state165_75_0 + shifted_state165_75_1 + shifted_state165_75_2 + shifted_state165_75_3 + shifted_state165_75_4 + shifted_state165_75_6 + shifted_state165_75_7 + shifted_state165_77_1 + shifted_state165_77_3 + shifted_state165_77_4 + shifted_state165_101_0 + shifted_state165_101_3 + shifted_state165_101_4 + shifted_state165_101_6 + shifted_state165_101_7 + shifted_state165_106_0 + shifted_state165_106_2 + shifted_state165_106_3 + shifted_state165_114_0 + shifted_state165_114_3 + shifted_state165_122_4 + shifted_state165_126_0 + shifted_state165_126_1 + shifted_state165_126_3 + shifted_state165_126_5 + shifted_state165_130_0 + shifted_state165_130_3 + shifted_state165_130_4 + shifted_state165_130_5 + shifted_state165_130_6 + shifted_state165_130_7 + shifted_state165_138_0 + shifted_state165_138_1 + shifted_state165_138_2 + shifted_state165_153_0 + shifted_state165_153_1 + shifted_state165_153_2 + shifted_state165_153_3 + shifted_state165_153_4 + shifted_state165_153_5 + shifted_state165_153_6 + shifted_state165_153_7 + shifted_state165_155_3 + shifted_state165_191_4 + shifted_state165_191_5 + shifted_state165_191_6 + shifted_state165_191_7 + shifted_state165_198_2 + shifted_state165_198_3 + shifted_state165_198_5 + shifted_state165_198_6 + shifted_state165_198_7);
      reservoir_sum_parallel[166] = (shifted_state166_0_2 + shifted_state166_0_3 + shifted_state166_0_4 + shifted_state166_0_5 + shifted_state166_0_6 + shifted_state166_0_7 + shifted_state166_3_0 + shifted_state166_3_2 + shifted_state166_3_4 + shifted_state166_16_4 + shifted_state166_16_6 + shifted_state166_16_7 + shifted_state166_17_2 + shifted_state166_17_3 + shifted_state166_17_5 + shifted_state166_17_6 + shifted_state166_17_7 + shifted_state166_26_0 + shifted_state166_26_1 + shifted_state166_26_2 + shifted_state166_26_5 + shifted_state166_26_6 + shifted_state166_26_7 + shifted_state166_29_3 + shifted_state166_29_5 + shifted_state166_29_6 + shifted_state166_29_7 + shifted_state166_32_0 + shifted_state166_32_1 + shifted_state166_32_2 + shifted_state166_32_3 + shifted_state166_32_5 + shifted_state166_32_6 + shifted_state166_32_7 + shifted_state166_38_0 + shifted_state166_38_1 + shifted_state166_38_2 + shifted_state166_38_6 + shifted_state166_45_3 + shifted_state166_45_4 + shifted_state166_45_5 + shifted_state166_46_1 + shifted_state166_46_2 + shifted_state166_46_3 + shifted_state166_46_5 + shifted_state166_46_6 + shifted_state166_46_7 + shifted_state166_50_1 + shifted_state166_50_5 + shifted_state166_50_6 + shifted_state166_50_7 + shifted_state166_74_2 + shifted_state166_74_4 + shifted_state166_95_3 + shifted_state166_95_4 + shifted_state166_95_5 + shifted_state166_95_6 + shifted_state166_95_7 + shifted_state166_98_0 + shifted_state166_98_1 + shifted_state166_98_3 + shifted_state166_111_2 + shifted_state166_111_5 + shifted_state166_111_6 + shifted_state166_111_7 + shifted_state166_116_2 + shifted_state166_116_5 + shifted_state166_116_6 + shifted_state166_116_7 + shifted_state166_121_3 + shifted_state166_121_5 + shifted_state166_121_6 + shifted_state166_121_7 + shifted_state166_123_0 + shifted_state166_123_2 + shifted_state166_123_4 + shifted_state166_127_0 + shifted_state166_127_1 + shifted_state166_127_4 + shifted_state166_127_5 + shifted_state166_127_6 + shifted_state166_127_7 + shifted_state166_158_1 + shifted_state166_158_3 + shifted_state166_158_4 + shifted_state166_158_5 + shifted_state166_158_6 + shifted_state166_158_7 + shifted_state166_168_0 + shifted_state166_170_5 + shifted_state166_170_6 + shifted_state166_170_7 + shifted_state166_187_0 + shifted_state166_187_3 + shifted_state166_187_4 + shifted_state166_187_5 + shifted_state166_187_6 + shifted_state166_187_7 + shifted_state166_191_0 + shifted_state166_191_2 + shifted_state166_191_4 + shifted_state166_191_5 + shifted_state166_192_0 + shifted_state166_192_4);
      reservoir_sum_parallel[167] = (shifted_state167_6_2 + shifted_state167_6_3 + shifted_state167_6_4 + shifted_state167_6_5 + shifted_state167_6_6 + shifted_state167_6_7 + shifted_state167_12_0 + shifted_state167_12_1 + shifted_state167_12_2 + shifted_state167_12_5 + shifted_state167_12_6 + shifted_state167_12_7 + shifted_state167_17_0 + shifted_state167_17_1 + shifted_state167_17_2 + shifted_state167_25_0 + shifted_state167_25_1 + shifted_state167_25_3 + shifted_state167_28_0 + shifted_state167_28_2 + shifted_state167_28_3 + shifted_state167_28_4 + shifted_state167_28_6 + shifted_state167_28_7 + shifted_state167_36_0 + shifted_state167_36_3 + shifted_state167_36_5 + shifted_state167_54_1 + shifted_state167_54_2 + shifted_state167_54_3 + shifted_state167_54_5 + shifted_state167_54_6 + shifted_state167_54_7 + shifted_state167_57_0 + shifted_state167_57_1 + shifted_state167_57_4 + shifted_state167_61_0 + shifted_state167_61_2 + shifted_state167_70_1 + shifted_state167_70_3 + shifted_state167_70_5 + shifted_state167_70_6 + shifted_state167_70_7 + shifted_state167_76_1 + shifted_state167_76_3 + shifted_state167_76_4 + shifted_state167_89_0 + shifted_state167_89_3 + shifted_state167_89_4 + shifted_state167_96_0 + shifted_state167_96_2 + shifted_state167_96_3 + shifted_state167_96_5 + shifted_state167_96_6 + shifted_state167_96_7 + shifted_state167_103_3 + shifted_state167_103_4 + shifted_state167_103_5 + shifted_state167_106_0 + shifted_state167_106_2 + shifted_state167_106_3 + shifted_state167_106_6 + shifted_state167_106_7 + shifted_state167_107_0 + shifted_state167_107_2 + shifted_state167_107_3 + shifted_state167_107_5 + shifted_state167_107_6 + shifted_state167_107_7 + shifted_state167_111_0 + shifted_state167_111_1 + shifted_state167_111_2 + shifted_state167_111_5 + shifted_state167_121_0 + shifted_state167_121_2 + shifted_state167_121_3 + shifted_state167_153_1 + shifted_state167_153_2 + shifted_state167_153_3 + shifted_state167_153_5 + shifted_state167_153_6 + shifted_state167_153_7 + shifted_state167_162_5 + shifted_state167_162_6 + shifted_state167_162_7 + shifted_state167_169_1 + shifted_state167_169_4 + shifted_state167_174_0 + shifted_state167_174_1 + shifted_state167_174_2 + shifted_state167_174_3 + shifted_state167_174_4 + shifted_state167_174_6 + shifted_state167_174_7 + shifted_state167_180_0 + shifted_state167_180_2 + shifted_state167_180_4 + shifted_state167_180_6 + shifted_state167_180_7 + shifted_state167_190_1 + shifted_state167_190_5 + shifted_state167_190_6 + shifted_state167_190_7 + shifted_state167_192_0 + shifted_state167_192_1 + shifted_state167_192_6 + shifted_state167_192_7 + shifted_state167_193_1 + shifted_state167_193_5 + shifted_state167_193_6 + shifted_state167_193_7);
      reservoir_sum_parallel[168] = (shifted_state168_7_0 + shifted_state168_7_1 + shifted_state168_11_0 + shifted_state168_11_2 + shifted_state168_19_1 + shifted_state168_19_2 + shifted_state168_19_3 + shifted_state168_20_0 + shifted_state168_20_2 + shifted_state168_20_3 + shifted_state168_20_4 + shifted_state168_20_5 + shifted_state168_20_6 + shifted_state168_20_7 + shifted_state168_28_0 + shifted_state168_28_1 + shifted_state168_28_4 + shifted_state168_31_2 + shifted_state168_31_5 + shifted_state168_31_6 + shifted_state168_31_7 + shifted_state168_39_1 + shifted_state168_39_2 + shifted_state168_39_3 + shifted_state168_39_6 + shifted_state168_39_7 + shifted_state168_41_0 + shifted_state168_41_1 + shifted_state168_41_3 + shifted_state168_41_4 + shifted_state168_41_5 + shifted_state168_41_6 + shifted_state168_41_7 + shifted_state168_56_0 + shifted_state168_56_1 + shifted_state168_56_4 + shifted_state168_63_0 + shifted_state168_63_3 + shifted_state168_63_4 + shifted_state168_63_6 + shifted_state168_63_7 + shifted_state168_68_1 + shifted_state168_68_3 + shifted_state168_93_0 + shifted_state168_93_5 + shifted_state168_93_6 + shifted_state168_93_7 + shifted_state168_140_1 + shifted_state168_141_2 + shifted_state168_141_3 + shifted_state168_141_4 + shifted_state168_141_5 + shifted_state168_141_6 + shifted_state168_141_7 + shifted_state168_142_2 + shifted_state168_142_5 + shifted_state168_177_0 + shifted_state168_177_1 + shifted_state168_180_0 + shifted_state168_180_2 + shifted_state168_180_3 + shifted_state168_180_5 + shifted_state168_180_6 + shifted_state168_180_7);
      reservoir_sum_parallel[169] = (shifted_state169_5_3 + shifted_state169_5_5 + shifted_state169_22_1 + shifted_state169_22_2 + shifted_state169_22_3 + shifted_state169_34_1 + shifted_state169_34_3 + shifted_state169_34_5 + shifted_state169_34_6 + shifted_state169_34_7 + shifted_state169_50_0 + shifted_state169_50_1 + shifted_state169_53_1 + shifted_state169_53_4 + shifted_state169_53_5 + shifted_state169_54_1 + shifted_state169_54_3 + shifted_state169_54_5 + shifted_state169_54_6 + shifted_state169_54_7 + shifted_state169_58_1 + shifted_state169_58_2 + shifted_state169_77_0 + shifted_state169_77_3 + shifted_state169_77_4 + shifted_state169_77_6 + shifted_state169_77_7 + shifted_state169_78_0 + shifted_state169_78_1 + shifted_state169_78_3 + shifted_state169_78_4 + shifted_state169_78_6 + shifted_state169_78_7 + shifted_state169_105_0 + shifted_state169_105_1 + shifted_state169_105_2 + shifted_state169_105_3 + shifted_state169_105_4 + shifted_state169_109_0 + shifted_state169_109_2 + shifted_state169_109_3 + shifted_state169_111_2 + shifted_state169_111_3 + shifted_state169_126_0 + shifted_state169_126_1 + shifted_state169_126_2 + shifted_state169_126_3 + shifted_state169_126_4 + shifted_state169_129_1 + shifted_state169_129_4 + shifted_state169_148_1 + shifted_state169_148_2 + shifted_state169_148_3 + shifted_state169_148_4 + shifted_state169_148_5 + shifted_state169_153_1 + shifted_state169_153_3 + shifted_state169_174_0 + shifted_state169_174_6);
      reservoir_sum_parallel[170] = (shifted_state170_12_0 + shifted_state170_12_1 + shifted_state170_12_5 + shifted_state170_12_6 + shifted_state170_12_7 + shifted_state170_22_0 + shifted_state170_22_1 + shifted_state170_22_2 + shifted_state170_22_4 + shifted_state170_22_5 + shifted_state170_22_6 + shifted_state170_22_7 + shifted_state170_34_1 + shifted_state170_34_2 + shifted_state170_34_5 + shifted_state170_66_0 + shifted_state170_66_2 + shifted_state170_66_3 + shifted_state170_66_4 + shifted_state170_66_6 + shifted_state170_70_2 + shifted_state170_70_3 + shifted_state170_70_5 + shifted_state170_70_6 + shifted_state170_70_7 + shifted_state170_81_0 + shifted_state170_81_3 + shifted_state170_81_4 + shifted_state170_97_5 + shifted_state170_97_6 + shifted_state170_97_7 + shifted_state170_98_0 + shifted_state170_98_1 + shifted_state170_98_2 + shifted_state170_98_4 + shifted_state170_98_5 + shifted_state170_98_6 + shifted_state170_98_7 + shifted_state170_104_1 + shifted_state170_104_2 + shifted_state170_104_3 + shifted_state170_104_4 + shifted_state170_106_2 + shifted_state170_106_4 + shifted_state170_106_5 + shifted_state170_118_2 + shifted_state170_118_5 + shifted_state170_118_6 + shifted_state170_118_7 + shifted_state170_124_0 + shifted_state170_124_1 + shifted_state170_133_0 + shifted_state170_133_2 + shifted_state170_140_1 + shifted_state170_140_4 + shifted_state170_140_5 + shifted_state170_140_6 + shifted_state170_140_7 + shifted_state170_162_1 + shifted_state170_162_4 + shifted_state170_162_5 + shifted_state170_162_6 + shifted_state170_162_7 + shifted_state170_172_0 + shifted_state170_172_1 + shifted_state170_172_2 + shifted_state170_172_3 + shifted_state170_173_1 + shifted_state170_173_3 + shifted_state170_173_4 + shifted_state170_173_5 + shifted_state170_173_6 + shifted_state170_173_7);
      reservoir_sum_parallel[171] = (shifted_state171_4_0 + shifted_state171_4_3 + shifted_state171_4_4 + shifted_state171_4_5 + shifted_state171_4_6 + shifted_state171_4_7 + shifted_state171_17_3 + shifted_state171_42_0 + shifted_state171_42_2 + shifted_state171_63_0 + shifted_state171_63_1 + shifted_state171_63_2 + shifted_state171_63_5 + shifted_state171_63_6 + shifted_state171_63_7 + shifted_state171_76_1 + shifted_state171_76_2 + shifted_state171_76_4 + shifted_state171_76_5 + shifted_state171_76_6 + shifted_state171_76_7 + shifted_state171_80_1 + shifted_state171_80_5 + shifted_state171_80_6 + shifted_state171_80_7 + shifted_state171_83_2 + shifted_state171_83_3 + shifted_state171_83_4 + shifted_state171_83_5 + shifted_state171_83_6 + shifted_state171_83_7 + shifted_state171_89_1 + shifted_state171_89_4 + shifted_state171_89_6 + shifted_state171_89_7 + shifted_state171_100_0 + shifted_state171_100_2 + shifted_state171_100_3 + shifted_state171_104_0 + shifted_state171_104_1 + shifted_state171_104_2 + shifted_state171_105_5 + shifted_state171_113_1 + shifted_state171_113_4 + shifted_state171_113_6 + shifted_state171_139_1 + shifted_state171_139_2 + shifted_state171_139_3 + shifted_state171_139_4 + shifted_state171_139_6 + shifted_state171_163_0 + shifted_state171_163_1 + shifted_state171_163_4 + shifted_state171_163_6 + shifted_state171_195_1 + shifted_state171_195_2 + shifted_state171_198_1 + shifted_state171_198_2 + shifted_state171_198_5 + shifted_state171_198_7);
      reservoir_sum_parallel[172] = (shifted_state172_5_0 + shifted_state172_5_1 + shifted_state172_5_2 + shifted_state172_5_4 + shifted_state172_5_5 + shifted_state172_5_6 + shifted_state172_5_7 + shifted_state172_8_2 + shifted_state172_8_4 + shifted_state172_8_5 + shifted_state172_8_6 + shifted_state172_8_7 + shifted_state172_20_2 + shifted_state172_20_5 + shifted_state172_20_6 + shifted_state172_20_7 + shifted_state172_28_0 + shifted_state172_28_1 + shifted_state172_32_2 + shifted_state172_32_3 + shifted_state172_32_4 + shifted_state172_32_5 + shifted_state172_35_0 + shifted_state172_54_0 + shifted_state172_54_1 + shifted_state172_54_2 + shifted_state172_54_3 + shifted_state172_54_4 + shifted_state172_66_3 + shifted_state172_66_4 + shifted_state172_66_5 + shifted_state172_66_6 + shifted_state172_66_7 + shifted_state172_72_1 + shifted_state172_72_5 + shifted_state172_72_6 + shifted_state172_72_7 + shifted_state172_89_0 + shifted_state172_89_2 + shifted_state172_89_3 + shifted_state172_89_4 + shifted_state172_89_5 + shifted_state172_89_6 + shifted_state172_89_7 + shifted_state172_112_1 + shifted_state172_112_5 + shifted_state172_119_1 + shifted_state172_119_3 + shifted_state172_119_5 + shifted_state172_128_0 + shifted_state172_128_1 + shifted_state172_128_3 + shifted_state172_132_0 + shifted_state172_132_2 + shifted_state172_132_3 + shifted_state172_132_5 + shifted_state172_134_1 + shifted_state172_134_3 + shifted_state172_134_5 + shifted_state172_134_6 + shifted_state172_134_7 + shifted_state172_164_0 + shifted_state172_164_3 + shifted_state172_164_5 + shifted_state172_164_6 + shifted_state172_164_7 + shifted_state172_167_2 + shifted_state172_175_0 + shifted_state172_175_1 + shifted_state172_175_2 + shifted_state172_175_3 + shifted_state172_175_4 + shifted_state172_191_1 + shifted_state172_194_0 + shifted_state172_194_2 + shifted_state172_194_3 + shifted_state172_194_4 + shifted_state172_194_6 + shifted_state172_194_7);
      reservoir_sum_parallel[173] = (shifted_state173_10_0 + shifted_state173_10_1 + shifted_state173_24_0 + shifted_state173_24_2 + shifted_state173_24_3 + shifted_state173_24_4 + shifted_state173_24_5 + shifted_state173_28_0 + shifted_state173_28_1 + shifted_state173_28_3 + shifted_state173_28_4 + shifted_state173_28_5 + shifted_state173_28_6 + shifted_state173_28_7 + shifted_state173_37_0 + shifted_state173_37_3 + shifted_state173_37_4 + shifted_state173_37_6 + shifted_state173_37_7 + shifted_state173_39_4 + shifted_state173_39_5 + shifted_state173_44_0 + shifted_state173_44_3 + shifted_state173_55_0 + shifted_state173_55_1 + shifted_state173_55_2 + shifted_state173_55_3 + shifted_state173_55_4 + shifted_state173_57_2 + shifted_state173_58_0 + shifted_state173_58_2 + shifted_state173_58_3 + shifted_state173_58_4 + shifted_state173_78_0 + shifted_state173_78_1 + shifted_state173_78_2 + shifted_state173_78_4 + shifted_state173_89_2 + shifted_state173_89_3 + shifted_state173_104_0 + shifted_state173_104_3 + shifted_state173_104_4 + shifted_state173_104_5 + shifted_state173_110_3 + shifted_state173_110_4 + shifted_state173_110_5 + shifted_state173_110_6 + shifted_state173_110_7 + shifted_state173_112_0 + shifted_state173_112_1 + shifted_state173_114_4 + shifted_state173_114_6 + shifted_state173_114_7 + shifted_state173_153_0 + shifted_state173_153_1 + shifted_state173_153_4 + shifted_state173_153_5);
      reservoir_sum_parallel[174] = (shifted_state174_10_0 + shifted_state174_10_3 + shifted_state174_14_1 + shifted_state174_14_2 + shifted_state174_18_0 + shifted_state174_18_1 + shifted_state174_31_1 + shifted_state174_31_3 + shifted_state174_31_5 + shifted_state174_32_0 + shifted_state174_57_1 + shifted_state174_57_3 + shifted_state174_57_4 + shifted_state174_57_6 + shifted_state174_57_7 + shifted_state174_63_0 + shifted_state174_63_1 + shifted_state174_63_2 + shifted_state174_63_5 + shifted_state174_63_6 + shifted_state174_63_7 + shifted_state174_64_3 + shifted_state174_64_4 + shifted_state174_79_0 + shifted_state174_79_1 + shifted_state174_88_1 + shifted_state174_88_2 + shifted_state174_88_3 + shifted_state174_113_2 + shifted_state174_113_3 + shifted_state174_113_5 + shifted_state174_113_6 + shifted_state174_113_7 + shifted_state174_115_2 + shifted_state174_115_3 + shifted_state174_115_5 + shifted_state174_144_2 + shifted_state174_144_3 + shifted_state174_145_0 + shifted_state174_145_1 + shifted_state174_145_2 + shifted_state174_145_3 + shifted_state174_148_1 + shifted_state174_148_2 + shifted_state174_148_4 + shifted_state174_151_3 + shifted_state174_151_4 + shifted_state174_151_5 + shifted_state174_151_6 + shifted_state174_151_7 + shifted_state174_154_1 + shifted_state174_154_4 + shifted_state174_154_5 + shifted_state174_154_6 + shifted_state174_154_7 + shifted_state174_155_2 + shifted_state174_155_4 + shifted_state174_155_5 + shifted_state174_163_0 + shifted_state174_163_5 + shifted_state174_166_0 + shifted_state174_166_1 + shifted_state174_166_3 + shifted_state174_166_4 + shifted_state174_170_0 + shifted_state174_170_2 + shifted_state174_170_3 + shifted_state174_170_4 + shifted_state174_170_5 + shifted_state174_170_6 + shifted_state174_170_7 + shifted_state174_171_1 + shifted_state174_171_2 + shifted_state174_171_3 + shifted_state174_192_2 + shifted_state174_192_3 + shifted_state174_192_4 + shifted_state174_192_5 + shifted_state174_192_6 + shifted_state174_192_7 + shifted_state174_198_0 + shifted_state174_198_1 + shifted_state174_198_2 + shifted_state174_198_5);
      reservoir_sum_parallel[175] = (shifted_state175_12_3 + shifted_state175_12_4 + shifted_state175_12_6 + shifted_state175_12_7 + shifted_state175_17_0 + shifted_state175_17_1 + shifted_state175_17_2 + shifted_state175_17_3 + shifted_state175_18_0 + shifted_state175_18_1 + shifted_state175_18_2 + shifted_state175_18_4 + shifted_state175_18_5 + shifted_state175_18_6 + shifted_state175_18_7 + shifted_state175_31_1 + shifted_state175_31_3 + shifted_state175_31_5 + shifted_state175_31_6 + shifted_state175_31_7 + shifted_state175_44_0 + shifted_state175_44_2 + shifted_state175_44_3 + shifted_state175_44_6 + shifted_state175_44_7 + shifted_state175_50_3 + shifted_state175_63_0 + shifted_state175_63_1 + shifted_state175_63_2 + shifted_state175_63_3 + shifted_state175_63_5 + shifted_state175_68_2 + shifted_state175_68_3 + shifted_state175_69_0 + shifted_state175_69_2 + shifted_state175_69_3 + shifted_state175_69_4 + shifted_state175_69_5 + shifted_state175_69_6 + shifted_state175_69_7 + shifted_state175_99_0 + shifted_state175_99_1 + shifted_state175_106_1 + shifted_state175_106_4 + shifted_state175_113_0 + shifted_state175_113_3 + shifted_state175_113_5 + shifted_state175_113_6 + shifted_state175_113_7 + shifted_state175_120_0 + shifted_state175_120_1 + shifted_state175_120_3 + shifted_state175_123_0 + shifted_state175_123_1 + shifted_state175_123_2 + shifted_state175_123_3 + shifted_state175_123_4 + shifted_state175_139_3 + shifted_state175_139_5 + shifted_state175_145_1 + shifted_state175_145_2 + shifted_state175_145_4 + shifted_state175_145_5 + shifted_state175_161_3 + shifted_state175_161_4 + shifted_state175_176_3 + shifted_state175_179_0 + shifted_state175_179_1 + shifted_state175_179_5 + shifted_state175_190_0 + shifted_state175_190_3 + shifted_state175_190_5 + shifted_state175_195_0 + shifted_state175_195_1 + shifted_state175_195_2 + shifted_state175_195_3);
      reservoir_sum_parallel[176] = (shifted_state176_28_3 + shifted_state176_28_4 + shifted_state176_28_5 + shifted_state176_28_6 + shifted_state176_28_7 + shifted_state176_38_1 + shifted_state176_38_4 + shifted_state176_70_0 + shifted_state176_70_1 + shifted_state176_70_3 + shifted_state176_70_5 + shifted_state176_70_6 + shifted_state176_70_7 + shifted_state176_79_1 + shifted_state176_79_4 + shifted_state176_94_1 + shifted_state176_94_2 + shifted_state176_94_3 + shifted_state176_94_4 + shifted_state176_94_5 + shifted_state176_94_6 + shifted_state176_94_7 + shifted_state176_110_0 + shifted_state176_110_1 + shifted_state176_110_3 + shifted_state176_115_0 + shifted_state176_115_2 + shifted_state176_115_5 + shifted_state176_130_0 + shifted_state176_130_1 + shifted_state176_130_2 + shifted_state176_130_5 + shifted_state176_133_4 + shifted_state176_140_0 + shifted_state176_140_1 + shifted_state176_140_3 + shifted_state176_140_4 + shifted_state176_144_3 + shifted_state176_144_4 + shifted_state176_144_5 + shifted_state176_144_6 + shifted_state176_144_7 + shifted_state176_146_1 + shifted_state176_146_4 + shifted_state176_146_6 + shifted_state176_148_0 + shifted_state176_148_1 + shifted_state176_148_3 + shifted_state176_148_5 + shifted_state176_148_6 + shifted_state176_148_7 + shifted_state176_173_0);
      reservoir_sum_parallel[177] = (shifted_state177_13_0 + shifted_state177_13_2 + shifted_state177_14_1 + shifted_state177_14_2 + shifted_state177_14_4 + shifted_state177_14_5 + shifted_state177_14_6 + shifted_state177_14_7 + shifted_state177_18_1 + shifted_state177_18_2 + shifted_state177_18_4 + shifted_state177_27_2 + shifted_state177_27_3 + shifted_state177_28_0 + shifted_state177_28_2 + shifted_state177_30_1 + shifted_state177_30_2 + shifted_state177_30_4 + shifted_state177_43_0 + shifted_state177_43_1 + shifted_state177_43_3 + shifted_state177_43_4 + shifted_state177_44_3 + shifted_state177_44_4 + shifted_state177_67_0 + shifted_state177_67_2 + shifted_state177_67_3 + shifted_state177_67_5 + shifted_state177_76_2 + shifted_state177_76_3 + shifted_state177_76_4 + shifted_state177_76_5 + shifted_state177_76_6 + shifted_state177_76_7 + shifted_state177_81_0 + shifted_state177_81_1 + shifted_state177_81_4 + shifted_state177_85_0 + shifted_state177_85_3 + shifted_state177_85_4 + shifted_state177_85_5 + shifted_state177_85_6 + shifted_state177_85_7 + shifted_state177_138_1 + shifted_state177_138_2 + shifted_state177_138_4 + shifted_state177_148_0 + shifted_state177_148_1 + shifted_state177_148_2 + shifted_state177_148_3 + shifted_state177_165_1 + shifted_state177_165_2 + shifted_state177_172_0 + shifted_state177_172_1 + shifted_state177_172_2 + shifted_state177_172_4 + shifted_state177_172_5 + shifted_state177_172_6 + shifted_state177_172_7 + shifted_state177_174_1 + shifted_state177_174_2 + shifted_state177_174_4 + shifted_state177_174_6 + shifted_state177_174_7 + shifted_state177_195_0 + shifted_state177_195_4 + shifted_state177_198_1 + shifted_state177_198_4 + shifted_state177_198_5 + shifted_state177_198_6 + shifted_state177_198_7);
      reservoir_sum_parallel[178] = (shifted_state178_19_2 + shifted_state178_19_4 + shifted_state178_19_5 + shifted_state178_19_6 + shifted_state178_19_7 + shifted_state178_21_0 + shifted_state178_21_1 + shifted_state178_21_4 + shifted_state178_21_6 + shifted_state178_21_7 + shifted_state178_60_0 + shifted_state178_60_1 + shifted_state178_60_2 + shifted_state178_60_5 + shifted_state178_60_6 + shifted_state178_60_7 + shifted_state178_61_0 + shifted_state178_61_4 + shifted_state178_82_0 + shifted_state178_82_1 + shifted_state178_82_2 + shifted_state178_82_5 + shifted_state178_82_6 + shifted_state178_82_7 + shifted_state178_87_0 + shifted_state178_87_1 + shifted_state178_87_2 + shifted_state178_87_4 + shifted_state178_87_6 + shifted_state178_87_7 + shifted_state178_92_1 + shifted_state178_92_2 + shifted_state178_92_3 + shifted_state178_93_3 + shifted_state178_93_4 + shifted_state178_93_6 + shifted_state178_93_7 + shifted_state178_110_0 + shifted_state178_110_2 + shifted_state178_110_3 + shifted_state178_133_0 + shifted_state178_133_1 + shifted_state178_133_4 + shifted_state178_133_5 + shifted_state178_133_6 + shifted_state178_133_7 + shifted_state178_136_1 + shifted_state178_138_4 + shifted_state178_138_5 + shifted_state178_138_6 + shifted_state178_138_7 + shifted_state178_144_0 + shifted_state178_144_1 + shifted_state178_144_3 + shifted_state178_144_4 + shifted_state178_144_5 + shifted_state178_164_1 + shifted_state178_164_2 + shifted_state178_164_3 + shifted_state178_164_4 + shifted_state178_164_5);
      reservoir_sum_parallel[179] = (shifted_state179_5_2 + shifted_state179_5_5 + shifted_state179_5_6 + shifted_state179_5_7 + shifted_state179_6_2 + shifted_state179_6_3 + shifted_state179_6_4 + shifted_state179_6_5 + shifted_state179_6_6 + shifted_state179_6_7 + shifted_state179_18_0 + shifted_state179_18_1 + shifted_state179_18_2 + shifted_state179_20_1 + shifted_state179_20_5 + shifted_state179_20_6 + shifted_state179_20_7 + shifted_state179_22_1 + shifted_state179_22_3 + shifted_state179_22_5 + shifted_state179_22_6 + shifted_state179_22_7 + shifted_state179_28_2 + shifted_state179_39_0 + shifted_state179_39_1 + shifted_state179_39_5 + shifted_state179_42_4 + shifted_state179_42_5 + shifted_state179_42_6 + shifted_state179_42_7 + shifted_state179_45_1 + shifted_state179_45_2 + shifted_state179_45_3 + shifted_state179_57_1 + shifted_state179_57_2 + shifted_state179_57_4 + shifted_state179_57_5 + shifted_state179_57_6 + shifted_state179_57_7 + shifted_state179_62_3 + shifted_state179_62_4 + shifted_state179_62_6 + shifted_state179_64_0 + shifted_state179_64_1 + shifted_state179_77_3 + shifted_state179_77_5 + shifted_state179_77_6 + shifted_state179_77_7 + shifted_state179_86_0 + shifted_state179_86_1 + shifted_state179_86_2 + shifted_state179_86_4 + shifted_state179_86_6 + shifted_state179_86_7 + shifted_state179_98_0 + shifted_state179_98_3 + shifted_state179_98_4 + shifted_state179_106_1 + shifted_state179_106_3 + shifted_state179_106_6 + shifted_state179_106_7 + shifted_state179_109_0 + shifted_state179_109_1 + shifted_state179_109_3 + shifted_state179_109_4 + shifted_state179_111_1 + shifted_state179_111_3 + shifted_state179_111_5 + shifted_state179_111_6 + shifted_state179_111_7 + shifted_state179_116_0 + shifted_state179_116_3 + shifted_state179_116_4 + shifted_state179_122_0 + shifted_state179_122_1 + shifted_state179_122_3 + shifted_state179_122_5 + shifted_state179_122_6 + shifted_state179_122_7 + shifted_state179_127_0 + shifted_state179_127_1 + shifted_state179_127_3 + shifted_state179_146_0 + shifted_state179_146_2 + shifted_state179_146_4 + shifted_state179_156_0 + shifted_state179_156_1 + shifted_state179_156_4 + shifted_state179_171_0 + shifted_state179_171_2 + shifted_state179_171_3 + shifted_state179_171_4 + shifted_state179_193_0 + shifted_state179_193_3 + shifted_state179_193_5 + shifted_state179_193_6 + shifted_state179_193_7);
      reservoir_sum_parallel[180] = (shifted_state180_0_1 + shifted_state180_0_2 + shifted_state180_0_3 + shifted_state180_0_4 + shifted_state180_0_5 + shifted_state180_0_6 + shifted_state180_0_7 + shifted_state180_3_0 + shifted_state180_3_1 + shifted_state180_3_4 + shifted_state180_18_0 + shifted_state180_18_2 + shifted_state180_18_3 + shifted_state180_18_4 + shifted_state180_18_5 + shifted_state180_18_6 + shifted_state180_18_7 + shifted_state180_32_0 + shifted_state180_32_1 + shifted_state180_32_2 + shifted_state180_33_0 + shifted_state180_33_1 + shifted_state180_33_4 + shifted_state180_38_0 + shifted_state180_38_2 + shifted_state180_38_5 + shifted_state180_39_0 + shifted_state180_39_1 + shifted_state180_39_3 + shifted_state180_39_4 + shifted_state180_39_5 + shifted_state180_39_6 + shifted_state180_39_7 + shifted_state180_41_0 + shifted_state180_41_1 + shifted_state180_41_2 + shifted_state180_41_3 + shifted_state180_41_4 + shifted_state180_42_0 + shifted_state180_42_5 + shifted_state180_42_6 + shifted_state180_42_7 + shifted_state180_49_1 + shifted_state180_49_2 + shifted_state180_49_3 + shifted_state180_49_4 + shifted_state180_49_5 + shifted_state180_49_6 + shifted_state180_49_7 + shifted_state180_66_0 + shifted_state180_66_1 + shifted_state180_66_3 + shifted_state180_66_4 + shifted_state180_66_5 + shifted_state180_66_6 + shifted_state180_66_7 + shifted_state180_73_0 + shifted_state180_73_4 + shifted_state180_73_6 + shifted_state180_73_7 + shifted_state180_76_0 + shifted_state180_76_1 + shifted_state180_76_2 + shifted_state180_76_4 + shifted_state180_76_6 + shifted_state180_76_7 + shifted_state180_77_1 + shifted_state180_77_2 + shifted_state180_77_3 + shifted_state180_77_5 + shifted_state180_77_6 + shifted_state180_77_7 + shifted_state180_86_1 + shifted_state180_95_0 + shifted_state180_95_3 + shifted_state180_95_5 + shifted_state180_95_6 + shifted_state180_95_7 + shifted_state180_99_0 + shifted_state180_99_1 + shifted_state180_99_2 + shifted_state180_99_4 + shifted_state180_106_2 + shifted_state180_112_1 + shifted_state180_112_4 + shifted_state180_112_5 + shifted_state180_112_6 + shifted_state180_112_7 + shifted_state180_113_1 + shifted_state180_113_2 + shifted_state180_113_4 + shifted_state180_121_0 + shifted_state180_121_1 + shifted_state180_121_3 + shifted_state180_127_2 + shifted_state180_127_3 + shifted_state180_127_5 + shifted_state180_127_6 + shifted_state180_127_7 + shifted_state180_143_2 + shifted_state180_143_5 + shifted_state180_143_6 + shifted_state180_143_7 + shifted_state180_145_0 + shifted_state180_145_2 + shifted_state180_145_3 + shifted_state180_147_0 + shifted_state180_147_3 + shifted_state180_147_4 + shifted_state180_160_0 + shifted_state180_160_5 + shifted_state180_161_1 + shifted_state180_161_3 + shifted_state180_161_4 + shifted_state180_164_0 + shifted_state180_164_2 + shifted_state180_164_5 + shifted_state180_164_6 + shifted_state180_164_7 + shifted_state180_190_0 + shifted_state180_190_1 + shifted_state180_190_2 + shifted_state180_190_5 + shifted_state180_192_0 + shifted_state180_192_1 + shifted_state180_192_2 + shifted_state180_192_3 + shifted_state180_192_4 + shifted_state180_192_5 + shifted_state180_192_6 + shifted_state180_192_7 + shifted_state180_193_0 + shifted_state180_193_2);
      reservoir_sum_parallel[181] = (shifted_state181_1_0 + shifted_state181_1_2 + shifted_state181_1_4 + shifted_state181_1_5 + shifted_state181_23_1 + shifted_state181_23_2 + shifted_state181_23_3 + shifted_state181_23_5 + shifted_state181_23_6 + shifted_state181_23_7 + shifted_state181_28_0 + shifted_state181_28_4 + shifted_state181_28_5 + shifted_state181_28_6 + shifted_state181_28_7 + shifted_state181_35_1 + shifted_state181_35_3 + shifted_state181_35_4 + shifted_state181_35_5 + shifted_state181_35_6 + shifted_state181_35_7 + shifted_state181_37_1 + shifted_state181_37_4 + shifted_state181_37_5 + shifted_state181_37_6 + shifted_state181_37_7 + shifted_state181_46_0 + shifted_state181_46_1 + shifted_state181_46_3 + shifted_state181_46_4 + shifted_state181_53_2 + shifted_state181_53_5 + shifted_state181_53_6 + shifted_state181_53_7 + shifted_state181_67_2 + shifted_state181_67_5 + shifted_state181_67_6 + shifted_state181_67_7 + shifted_state181_73_1 + shifted_state181_73_4 + shifted_state181_74_0 + shifted_state181_74_1 + shifted_state181_74_2 + shifted_state181_74_5 + shifted_state181_74_6 + shifted_state181_74_7 + shifted_state181_80_2 + shifted_state181_80_3 + shifted_state181_80_5 + shifted_state181_80_6 + shifted_state181_80_7 + shifted_state181_85_0 + shifted_state181_85_1 + shifted_state181_85_3 + shifted_state181_92_0 + shifted_state181_92_2 + shifted_state181_92_4 + shifted_state181_92_6 + shifted_state181_92_7 + shifted_state181_98_0 + shifted_state181_104_3 + shifted_state181_104_4 + shifted_state181_104_5 + shifted_state181_137_0 + shifted_state181_137_2 + shifted_state181_137_3 + shifted_state181_137_5 + shifted_state181_144_2 + shifted_state181_144_3 + shifted_state181_144_5 + shifted_state181_150_0 + shifted_state181_150_2 + shifted_state181_150_3 + shifted_state181_150_5 + shifted_state181_150_6 + shifted_state181_150_7 + shifted_state181_151_1 + shifted_state181_151_2 + shifted_state181_151_3 + shifted_state181_151_5 + shifted_state181_151_6 + shifted_state181_151_7 + shifted_state181_168_1 + shifted_state181_168_2 + shifted_state181_168_4 + shifted_state181_168_5 + shifted_state181_168_6 + shifted_state181_168_7 + shifted_state181_175_1 + shifted_state181_175_3 + shifted_state181_190_0 + shifted_state181_190_1 + shifted_state181_190_2 + shifted_state181_190_4 + shifted_state181_190_5 + shifted_state181_190_6 + shifted_state181_190_7);
      reservoir_sum_parallel[182] = (shifted_state182_26_3 + shifted_state182_27_0 + shifted_state182_27_6 + shifted_state182_27_7 + shifted_state182_36_0 + shifted_state182_36_4 + shifted_state182_36_5 + shifted_state182_36_6 + shifted_state182_36_7 + shifted_state182_48_0 + shifted_state182_48_2 + shifted_state182_48_3 + shifted_state182_48_4 + shifted_state182_52_2 + shifted_state182_52_4 + shifted_state182_52_5 + shifted_state182_64_1 + shifted_state182_64_2 + shifted_state182_64_3 + shifted_state182_64_5 + shifted_state182_65_1 + shifted_state182_65_4 + shifted_state182_65_5 + shifted_state182_93_1 + shifted_state182_93_4 + shifted_state182_99_0 + shifted_state182_99_3 + shifted_state182_99_4 + shifted_state182_99_5 + shifted_state182_99_6 + shifted_state182_99_7 + shifted_state182_132_2 + shifted_state182_132_3 + shifted_state182_132_5 + shifted_state182_145_0 + shifted_state182_145_2 + shifted_state182_166_2 + shifted_state182_166_4 + shifted_state182_175_1 + shifted_state182_175_3 + shifted_state182_175_5 + shifted_state182_175_6 + shifted_state182_175_7 + shifted_state182_178_2 + shifted_state182_178_3 + shifted_state182_178_4 + shifted_state182_178_5 + shifted_state182_185_2 + shifted_state182_185_3 + shifted_state182_185_5 + shifted_state182_185_6 + shifted_state182_185_7 + shifted_state182_186_1 + shifted_state182_186_3 + shifted_state182_186_4 + shifted_state182_187_3 + shifted_state182_187_5 + shifted_state182_187_6 + shifted_state182_187_7 + shifted_state182_197_1 + shifted_state182_197_3 + shifted_state182_197_6 + shifted_state182_197_7);
      reservoir_sum_parallel[183] = (shifted_state183_10_1 + shifted_state183_10_2 + shifted_state183_10_3 + shifted_state183_25_2 + shifted_state183_25_3 + shifted_state183_25_5 + shifted_state183_37_1 + shifted_state183_37_3 + shifted_state183_37_6 + shifted_state183_37_7 + shifted_state183_44_2 + shifted_state183_44_3 + shifted_state183_52_3 + shifted_state183_52_4 + shifted_state183_52_5 + shifted_state183_52_6 + shifted_state183_52_7 + shifted_state183_58_3 + shifted_state183_64_2 + shifted_state183_64_5 + shifted_state183_95_0 + shifted_state183_95_2 + shifted_state183_95_3 + shifted_state183_95_4 + shifted_state183_95_6 + shifted_state183_95_7 + shifted_state183_97_1 + shifted_state183_97_3 + shifted_state183_97_5 + shifted_state183_110_1 + shifted_state183_110_3 + shifted_state183_126_2 + shifted_state183_126_4 + shifted_state183_126_5 + shifted_state183_126_6 + shifted_state183_126_7 + shifted_state183_131_0 + shifted_state183_131_1 + shifted_state183_131_2 + shifted_state183_131_3 + shifted_state183_140_1 + shifted_state183_140_4 + shifted_state183_140_5 + shifted_state183_140_6 + shifted_state183_140_7 + shifted_state183_144_1 + shifted_state183_144_3 + shifted_state183_144_4 + shifted_state183_161_1 + shifted_state183_161_2 + shifted_state183_161_4 + shifted_state183_161_5 + shifted_state183_161_6 + shifted_state183_161_7 + shifted_state183_165_0 + shifted_state183_165_1 + shifted_state183_165_3 + shifted_state183_165_4 + shifted_state183_165_5 + shifted_state183_165_6 + shifted_state183_165_7 + shifted_state183_167_2 + shifted_state183_167_3 + shifted_state183_195_2 + shifted_state183_195_3);
      reservoir_sum_parallel[184] = (shifted_state184_2_1 + shifted_state184_2_3 + shifted_state184_2_6 + shifted_state184_2_7 + shifted_state184_28_0 + shifted_state184_28_2 + shifted_state184_28_3 + shifted_state184_28_4 + shifted_state184_31_1 + shifted_state184_31_2 + shifted_state184_31_5 + shifted_state184_31_6 + shifted_state184_31_7 + shifted_state184_34_4 + shifted_state184_35_0 + shifted_state184_35_1 + shifted_state184_35_5 + shifted_state184_35_6 + shifted_state184_35_7 + shifted_state184_37_0 + shifted_state184_37_4 + shifted_state184_37_6 + shifted_state184_37_7 + shifted_state184_39_2 + shifted_state184_39_3 + shifted_state184_39_4 + shifted_state184_42_0 + shifted_state184_42_1 + shifted_state184_42_3 + shifted_state184_42_4 + shifted_state184_42_6 + shifted_state184_42_7 + shifted_state184_45_0 + shifted_state184_46_0 + shifted_state184_46_2 + shifted_state184_46_3 + shifted_state184_50_3 + shifted_state184_52_1 + shifted_state184_52_2 + shifted_state184_52_4 + shifted_state184_52_5 + shifted_state184_52_6 + shifted_state184_52_7 + shifted_state184_70_1 + shifted_state184_70_2 + shifted_state184_70_5 + shifted_state184_70_6 + shifted_state184_70_7 + shifted_state184_71_2 + shifted_state184_71_5 + shifted_state184_71_6 + shifted_state184_71_7 + shifted_state184_83_0 + shifted_state184_83_1 + shifted_state184_83_2 + shifted_state184_83_4 + shifted_state184_101_0 + shifted_state184_101_1 + shifted_state184_101_2 + shifted_state184_101_3 + shifted_state184_101_5 + shifted_state184_101_6 + shifted_state184_101_7 + shifted_state184_114_0 + shifted_state184_114_1 + shifted_state184_114_3 + shifted_state184_114_4 + shifted_state184_117_0 + shifted_state184_117_1 + shifted_state184_117_3 + shifted_state184_117_4 + shifted_state184_117_6 + shifted_state184_117_7 + shifted_state184_134_1 + shifted_state184_134_3 + shifted_state184_134_6 + shifted_state184_134_7 + shifted_state184_140_0 + shifted_state184_140_1 + shifted_state184_140_2 + shifted_state184_165_0 + shifted_state184_165_3 + shifted_state184_165_6 + shifted_state184_165_7 + shifted_state184_171_1 + shifted_state184_171_2 + shifted_state184_171_4 + shifted_state184_192_0 + shifted_state184_192_1 + shifted_state184_192_3 + shifted_state184_192_5 + shifted_state184_192_6 + shifted_state184_192_7 + shifted_state184_193_1 + shifted_state184_193_4 + shifted_state184_193_5);
      reservoir_sum_parallel[185] = (shifted_state185_2_0 + shifted_state185_2_1 + shifted_state185_2_5 + shifted_state185_2_6 + shifted_state185_2_7 + shifted_state185_6_0 + shifted_state185_6_2 + shifted_state185_6_3 + shifted_state185_6_4 + shifted_state185_6_6 + shifted_state185_6_7 + shifted_state185_11_0 + shifted_state185_11_1 + shifted_state185_11_4 + shifted_state185_15_4 + shifted_state185_15_6 + shifted_state185_15_7 + shifted_state185_46_3 + shifted_state185_46_5 + shifted_state185_47_1 + shifted_state185_49_2 + shifted_state185_49_3 + shifted_state185_49_5 + shifted_state185_49_6 + shifted_state185_49_7 + shifted_state185_50_1 + shifted_state185_50_4 + shifted_state185_50_6 + shifted_state185_50_7 + shifted_state185_69_0 + shifted_state185_69_3 + shifted_state185_69_4 + shifted_state185_87_0 + shifted_state185_87_1 + shifted_state185_87_2 + shifted_state185_87_4 + shifted_state185_87_5 + shifted_state185_87_6 + shifted_state185_87_7 + shifted_state185_93_0 + shifted_state185_93_1 + shifted_state185_93_2 + shifted_state185_97_0 + shifted_state185_97_5 + shifted_state185_97_6 + shifted_state185_97_7 + shifted_state185_115_1 + shifted_state185_115_4 + shifted_state185_116_0 + shifted_state185_116_1 + shifted_state185_133_1 + shifted_state185_133_3 + shifted_state185_133_4 + shifted_state185_160_1 + shifted_state185_160_3 + shifted_state185_169_1 + shifted_state185_169_4 + shifted_state185_169_5 + shifted_state185_169_6 + shifted_state185_169_7 + shifted_state185_185_1 + shifted_state185_185_3 + shifted_state185_185_4);
      reservoir_sum_parallel[186] = (shifted_state186_8_0 + shifted_state186_8_1 + shifted_state186_8_2 + shifted_state186_8_3 + shifted_state186_10_0 + shifted_state186_10_1 + shifted_state186_10_2 + shifted_state186_10_3 + shifted_state186_10_5 + shifted_state186_10_6 + shifted_state186_10_7 + shifted_state186_14_4 + shifted_state186_14_6 + shifted_state186_14_7 + shifted_state186_39_1 + shifted_state186_39_3 + shifted_state186_45_0 + shifted_state186_45_1 + shifted_state186_45_2 + shifted_state186_45_3 + shifted_state186_51_0 + shifted_state186_51_2 + shifted_state186_51_3 + shifted_state186_63_0 + shifted_state186_63_3 + shifted_state186_63_4 + shifted_state186_63_6 + shifted_state186_63_7 + shifted_state186_73_0 + shifted_state186_73_1 + shifted_state186_73_2 + shifted_state186_73_3 + shifted_state186_73_4 + shifted_state186_83_0 + shifted_state186_83_3 + shifted_state186_83_4 + shifted_state186_83_6 + shifted_state186_83_7 + shifted_state186_85_0 + shifted_state186_85_6 + shifted_state186_86_3 + shifted_state186_86_6 + shifted_state186_86_7 + shifted_state186_88_0 + shifted_state186_88_1 + shifted_state186_88_2 + shifted_state186_88_4 + shifted_state186_110_0 + shifted_state186_110_2 + shifted_state186_110_3 + shifted_state186_110_5 + shifted_state186_110_6 + shifted_state186_110_7 + shifted_state186_125_1 + shifted_state186_125_2 + shifted_state186_125_3 + shifted_state186_125_6 + shifted_state186_125_7 + shifted_state186_127_1 + shifted_state186_133_5 + shifted_state186_147_0 + shifted_state186_147_1 + shifted_state186_147_2 + shifted_state186_147_3 + shifted_state186_147_4 + shifted_state186_153_1 + shifted_state186_153_3 + shifted_state186_153_6 + shifted_state186_156_0 + shifted_state186_156_1 + shifted_state186_156_2 + shifted_state186_156_3 + shifted_state186_163_0 + shifted_state186_163_1 + shifted_state186_163_2);
      reservoir_sum_parallel[187] = (shifted_state187_11_1 + shifted_state187_11_2 + shifted_state187_11_4 + shifted_state187_11_5 + shifted_state187_11_6 + shifted_state187_11_7 + shifted_state187_12_0 + shifted_state187_12_2 + shifted_state187_12_3 + shifted_state187_12_5 + shifted_state187_20_1 + shifted_state187_20_2 + shifted_state187_40_0 + shifted_state187_40_3 + shifted_state187_40_5 + shifted_state187_40_6 + shifted_state187_40_7 + shifted_state187_41_0 + shifted_state187_41_3 + shifted_state187_49_1 + shifted_state187_49_5 + shifted_state187_49_6 + shifted_state187_49_7 + shifted_state187_58_3 + shifted_state187_60_1 + shifted_state187_60_2 + shifted_state187_60_4 + shifted_state187_60_5 + shifted_state187_60_6 + shifted_state187_60_7 + shifted_state187_62_0 + shifted_state187_62_3 + shifted_state187_86_2 + shifted_state187_86_4 + shifted_state187_86_5 + shifted_state187_86_6 + shifted_state187_86_7 + shifted_state187_97_0 + shifted_state187_97_2 + shifted_state187_97_3 + shifted_state187_97_4 + shifted_state187_97_5 + shifted_state187_97_6 + shifted_state187_97_7 + shifted_state187_100_0 + shifted_state187_100_2 + shifted_state187_100_3 + shifted_state187_100_5 + shifted_state187_100_6 + shifted_state187_100_7 + shifted_state187_105_0 + shifted_state187_105_1 + shifted_state187_105_2 + shifted_state187_105_4 + shifted_state187_105_5 + shifted_state187_105_6 + shifted_state187_105_7 + shifted_state187_111_1 + shifted_state187_137_0 + shifted_state187_137_1 + shifted_state187_137_3 + shifted_state187_137_4 + shifted_state187_137_6 + shifted_state187_137_7 + shifted_state187_140_0 + shifted_state187_140_1 + shifted_state187_140_2 + shifted_state187_140_3 + shifted_state187_140_5 + shifted_state187_140_6 + shifted_state187_140_7 + shifted_state187_147_1 + shifted_state187_147_4 + shifted_state187_147_6 + shifted_state187_147_7 + shifted_state187_150_0 + shifted_state187_150_1 + shifted_state187_150_3 + shifted_state187_150_4 + shifted_state187_150_5 + shifted_state187_150_6 + shifted_state187_150_7 + shifted_state187_171_2 + shifted_state187_171_3 + shifted_state187_171_4 + shifted_state187_183_0 + shifted_state187_183_1 + shifted_state187_183_2 + shifted_state187_183_4 + shifted_state187_183_5 + shifted_state187_183_6 + shifted_state187_183_7 + shifted_state187_188_2 + shifted_state187_188_3 + shifted_state187_188_5 + shifted_state187_188_6 + shifted_state187_188_7);
      reservoir_sum_parallel[188] = (shifted_state188_4_1 + shifted_state188_4_2 + shifted_state188_4_4 + shifted_state188_4_5 + shifted_state188_4_6 + shifted_state188_4_7 + shifted_state188_5_2 + shifted_state188_5_3 + shifted_state188_5_5 + shifted_state188_5_6 + shifted_state188_5_7 + shifted_state188_18_0 + shifted_state188_18_1 + shifted_state188_18_2 + shifted_state188_18_3 + shifted_state188_18_4 + shifted_state188_18_5 + shifted_state188_18_6 + shifted_state188_18_7 + shifted_state188_33_1 + shifted_state188_33_2 + shifted_state188_33_5 + shifted_state188_33_6 + shifted_state188_33_7 + shifted_state188_42_0 + shifted_state188_42_1 + shifted_state188_42_2 + shifted_state188_42_4 + shifted_state188_42_6 + shifted_state188_42_7 + shifted_state188_44_2 + shifted_state188_44_4 + shifted_state188_44_6 + shifted_state188_44_7 + shifted_state188_45_1 + shifted_state188_45_2 + shifted_state188_63_1 + shifted_state188_63_2 + shifted_state188_63_3 + shifted_state188_63_5 + shifted_state188_63_6 + shifted_state188_63_7 + shifted_state188_89_2 + shifted_state188_89_5 + shifted_state188_89_6 + shifted_state188_89_7 + shifted_state188_100_5 + shifted_state188_104_2 + shifted_state188_104_5 + shifted_state188_104_6 + shifted_state188_104_7 + shifted_state188_106_1 + shifted_state188_106_2 + shifted_state188_106_3 + shifted_state188_106_4 + shifted_state188_116_1 + shifted_state188_116_2 + shifted_state188_116_3 + shifted_state188_116_4 + shifted_state188_116_5 + shifted_state188_116_6 + shifted_state188_116_7 + shifted_state188_117_0 + shifted_state188_117_3 + shifted_state188_117_4 + shifted_state188_117_6 + shifted_state188_117_7 + shifted_state188_127_0 + shifted_state188_127_3 + shifted_state188_127_4 + shifted_state188_127_5 + shifted_state188_127_6 + shifted_state188_127_7 + shifted_state188_130_4 + shifted_state188_130_6 + shifted_state188_130_7 + shifted_state188_142_1 + shifted_state188_142_2 + shifted_state188_142_3 + shifted_state188_142_5 + shifted_state188_142_6 + shifted_state188_142_7 + shifted_state188_150_0 + shifted_state188_150_2 + shifted_state188_150_3 + shifted_state188_150_4 + shifted_state188_155_1 + shifted_state188_155_2 + shifted_state188_186_0 + shifted_state188_186_2 + shifted_state188_186_3 + shifted_state188_186_4 + shifted_state188_186_6 + shifted_state188_186_7 + shifted_state188_192_0 + shifted_state188_192_2 + shifted_state188_192_4 + shifted_state188_192_5 + shifted_state188_192_6 + shifted_state188_192_7 + shifted_state188_195_0 + shifted_state188_195_5 + shifted_state188_197_2 + shifted_state188_197_3 + shifted_state188_197_4 + shifted_state188_197_6 + shifted_state188_197_7);
      reservoir_sum_parallel[189] = (shifted_state189_14_0 + shifted_state189_14_1 + shifted_state189_14_2 + shifted_state189_21_0 + shifted_state189_21_5 + shifted_state189_36_0 + shifted_state189_36_1 + shifted_state189_36_2 + shifted_state189_36_3 + shifted_state189_36_4 + shifted_state189_36_5 + shifted_state189_36_6 + shifted_state189_36_7 + shifted_state189_39_1 + shifted_state189_39_2 + shifted_state189_39_3 + shifted_state189_41_0 + shifted_state189_41_2 + shifted_state189_41_4 + shifted_state189_41_5 + shifted_state189_41_6 + shifted_state189_41_7 + shifted_state189_48_2 + shifted_state189_48_3 + shifted_state189_67_1 + shifted_state189_67_2 + shifted_state189_67_3 + shifted_state189_67_4 + shifted_state189_72_3 + shifted_state189_72_4 + shifted_state189_72_5 + shifted_state189_72_6 + shifted_state189_72_7 + shifted_state189_78_3 + shifted_state189_78_4 + shifted_state189_78_5 + shifted_state189_78_6 + shifted_state189_78_7 + shifted_state189_95_0 + shifted_state189_95_1 + shifted_state189_95_2 + shifted_state189_95_3 + shifted_state189_127_1 + shifted_state189_127_2 + shifted_state189_127_4 + shifted_state189_127_5 + shifted_state189_127_6 + shifted_state189_127_7 + shifted_state189_130_0 + shifted_state189_130_1 + shifted_state189_130_2 + shifted_state189_130_3 + shifted_state189_141_0 + shifted_state189_141_2 + shifted_state189_141_6 + shifted_state189_141_7 + shifted_state189_150_0 + shifted_state189_150_1 + shifted_state189_150_2 + shifted_state189_161_1 + shifted_state189_161_2 + shifted_state189_161_3 + shifted_state189_161_5 + shifted_state189_161_6 + shifted_state189_161_7 + shifted_state189_179_1 + shifted_state189_189_0 + shifted_state189_189_3 + shifted_state189_194_1 + shifted_state189_194_3 + shifted_state189_194_5 + shifted_state189_194_6 + shifted_state189_194_7 + shifted_state189_196_0 + shifted_state189_196_2 + shifted_state189_196_3 + shifted_state189_196_4 + shifted_state189_196_6 + shifted_state189_196_7);
      reservoir_sum_parallel[190] = (shifted_state190_11_0 + shifted_state190_11_2 + shifted_state190_11_3 + shifted_state190_11_4 + shifted_state190_11_5 + shifted_state190_11_6 + shifted_state190_11_7 + shifted_state190_15_3 + shifted_state190_15_5 + shifted_state190_15_6 + shifted_state190_15_7 + shifted_state190_21_0 + shifted_state190_21_1 + shifted_state190_21_4 + shifted_state190_21_5 + shifted_state190_62_2 + shifted_state190_65_0 + shifted_state190_65_1 + shifted_state190_65_2 + shifted_state190_65_5 + shifted_state190_65_6 + shifted_state190_65_7 + shifted_state190_66_1 + shifted_state190_66_3 + shifted_state190_66_4 + shifted_state190_80_0 + shifted_state190_80_1 + shifted_state190_80_2 + shifted_state190_80_4 + shifted_state190_80_5 + shifted_state190_91_0 + shifted_state190_91_2 + shifted_state190_91_3 + shifted_state190_91_4 + shifted_state190_91_6 + shifted_state190_91_7 + shifted_state190_97_0 + shifted_state190_97_3 + shifted_state190_97_4 + shifted_state190_107_1 + shifted_state190_107_3 + shifted_state190_107_5 + shifted_state190_107_6 + shifted_state190_107_7 + shifted_state190_109_2 + shifted_state190_109_3 + shifted_state190_109_6 + shifted_state190_109_7 + shifted_state190_160_0 + shifted_state190_160_2 + shifted_state190_163_3 + shifted_state190_172_0 + shifted_state190_172_1 + shifted_state190_172_2 + shifted_state190_172_3 + shifted_state190_172_5 + shifted_state190_175_0 + shifted_state190_175_5 + shifted_state190_175_6 + shifted_state190_175_7 + shifted_state190_189_1 + shifted_state190_189_2 + shifted_state190_189_3 + shifted_state190_189_5 + shifted_state190_189_6 + shifted_state190_189_7 + shifted_state190_194_4 + shifted_state190_199_0 + shifted_state190_199_1 + shifted_state190_199_3 + shifted_state190_199_5 + shifted_state190_199_6 + shifted_state190_199_7);
      reservoir_sum_parallel[191] = (shifted_state191_1_1 + shifted_state191_1_2 + shifted_state191_1_6 + shifted_state191_4_0 + shifted_state191_6_0 + shifted_state191_6_1 + shifted_state191_6_2 + shifted_state191_6_3 + shifted_state191_13_0 + shifted_state191_13_1 + shifted_state191_13_3 + shifted_state191_13_5 + shifted_state191_13_6 + shifted_state191_13_7 + shifted_state191_26_2 + shifted_state191_26_3 + shifted_state191_26_4 + shifted_state191_30_0 + shifted_state191_30_2 + shifted_state191_30_3 + shifted_state191_30_4 + shifted_state191_30_5 + shifted_state191_30_6 + shifted_state191_30_7 + shifted_state191_43_4 + shifted_state191_43_5 + shifted_state191_43_6 + shifted_state191_43_7 + shifted_state191_45_0 + shifted_state191_45_1 + shifted_state191_45_4 + shifted_state191_45_5 + shifted_state191_45_6 + shifted_state191_45_7 + shifted_state191_56_1 + shifted_state191_59_1 + shifted_state191_59_2 + shifted_state191_59_3 + shifted_state191_59_4 + shifted_state191_59_5 + shifted_state191_59_6 + shifted_state191_59_7 + shifted_state191_69_0 + shifted_state191_69_1 + shifted_state191_69_3 + shifted_state191_84_0 + shifted_state191_84_1 + shifted_state191_84_2 + shifted_state191_98_0 + shifted_state191_98_2 + shifted_state191_98_3 + shifted_state191_98_4 + shifted_state191_98_5 + shifted_state191_106_3 + shifted_state191_106_5 + shifted_state191_106_6 + shifted_state191_106_7 + shifted_state191_132_0 + shifted_state191_132_1 + shifted_state191_132_2 + shifted_state191_132_4 + shifted_state191_147_0 + shifted_state191_147_4 + shifted_state191_147_5 + shifted_state191_168_0 + shifted_state191_169_4 + shifted_state191_174_2 + shifted_state191_174_4 + shifted_state191_174_6 + shifted_state191_174_7 + shifted_state191_179_1 + shifted_state191_179_2 + shifted_state191_179_3 + shifted_state191_179_5 + shifted_state191_187_0 + shifted_state191_187_1 + shifted_state191_187_2 + shifted_state191_187_3 + shifted_state191_187_4 + shifted_state191_187_5 + shifted_state191_187_6 + shifted_state191_187_7 + shifted_state191_194_0 + shifted_state191_194_2 + shifted_state191_194_3 + shifted_state191_194_6 + shifted_state191_194_7 + shifted_state191_197_1 + shifted_state191_197_3 + shifted_state191_197_4);
      reservoir_sum_parallel[192] = (shifted_state192_1_0 + shifted_state192_1_1 + shifted_state192_1_2 + shifted_state192_1_3 + shifted_state192_1_4 + shifted_state192_1_5 + shifted_state192_1_6 + shifted_state192_1_7 + shifted_state192_19_0 + shifted_state192_19_2 + shifted_state192_19_3 + shifted_state192_19_5 + shifted_state192_19_6 + shifted_state192_19_7 + shifted_state192_22_0 + shifted_state192_22_2 + shifted_state192_22_4 + shifted_state192_22_5 + shifted_state192_22_6 + shifted_state192_22_7 + shifted_state192_24_0 + shifted_state192_24_1 + shifted_state192_24_2 + shifted_state192_24_4 + shifted_state192_24_5 + shifted_state192_24_6 + shifted_state192_24_7 + shifted_state192_31_0 + shifted_state192_31_4 + shifted_state192_31_5 + shifted_state192_44_0 + shifted_state192_44_2 + shifted_state192_54_1 + shifted_state192_54_4 + shifted_state192_63_0 + shifted_state192_63_3 + shifted_state192_63_5 + shifted_state192_63_6 + shifted_state192_63_7 + shifted_state192_77_3 + shifted_state192_77_4 + shifted_state192_77_5 + shifted_state192_77_6 + shifted_state192_77_7 + shifted_state192_81_0 + shifted_state192_81_1 + shifted_state192_81_3 + shifted_state192_81_4 + shifted_state192_81_5 + shifted_state192_81_6 + shifted_state192_81_7 + shifted_state192_93_0 + shifted_state192_93_1 + shifted_state192_93_3 + shifted_state192_93_5 + shifted_state192_94_1 + shifted_state192_94_2 + shifted_state192_95_4 + shifted_state192_95_5 + shifted_state192_95_6 + shifted_state192_95_7 + shifted_state192_96_2 + shifted_state192_96_4 + shifted_state192_96_5 + shifted_state192_96_6 + shifted_state192_96_7 + shifted_state192_103_1 + shifted_state192_103_4 + shifted_state192_103_6 + shifted_state192_103_7 + shifted_state192_112_2 + shifted_state192_112_3 + shifted_state192_112_5 + shifted_state192_112_6 + shifted_state192_112_7 + shifted_state192_114_2 + shifted_state192_114_3 + shifted_state192_116_0 + shifted_state192_116_2 + shifted_state192_116_3 + shifted_state192_116_4 + shifted_state192_118_0 + shifted_state192_118_1 + shifted_state192_118_2 + shifted_state192_118_4 + shifted_state192_118_5 + shifted_state192_118_6 + shifted_state192_118_7 + shifted_state192_123_0 + shifted_state192_123_1 + shifted_state192_123_3 + shifted_state192_123_4 + shifted_state192_123_5 + shifted_state192_123_6 + shifted_state192_123_7 + shifted_state192_136_1 + shifted_state192_136_2 + shifted_state192_136_4 + shifted_state192_136_5 + shifted_state192_136_6 + shifted_state192_136_7 + shifted_state192_161_0 + shifted_state192_161_1 + shifted_state192_161_4 + shifted_state192_161_5 + shifted_state192_161_6 + shifted_state192_161_7 + shifted_state192_166_2 + shifted_state192_166_4 + shifted_state192_166_6 + shifted_state192_166_7);
      reservoir_sum_parallel[193] = (shifted_state193_1_2 + shifted_state193_4_0 + shifted_state193_16_0 + shifted_state193_16_4 + shifted_state193_39_1 + shifted_state193_39_4 + shifted_state193_39_5 + shifted_state193_41_1 + shifted_state193_41_2 + shifted_state193_41_3 + shifted_state193_41_4 + shifted_state193_41_5 + shifted_state193_41_6 + shifted_state193_41_7 + shifted_state193_50_1 + shifted_state193_51_0 + shifted_state193_51_1 + shifted_state193_51_2 + shifted_state193_51_3 + shifted_state193_51_5 + shifted_state193_67_0 + shifted_state193_67_1 + shifted_state193_67_2 + shifted_state193_67_4 + shifted_state193_67_6 + shifted_state193_67_7 + shifted_state193_84_2 + shifted_state193_84_3 + shifted_state193_86_0 + shifted_state193_86_4 + shifted_state193_89_0 + shifted_state193_89_2 + shifted_state193_90_1 + shifted_state193_90_2 + shifted_state193_90_6 + shifted_state193_90_7 + shifted_state193_100_2 + shifted_state193_100_3 + shifted_state193_100_4 + shifted_state193_101_2 + shifted_state193_101_3 + shifted_state193_101_4 + shifted_state193_101_5 + shifted_state193_101_6 + shifted_state193_101_7 + shifted_state193_102_0 + shifted_state193_102_1 + shifted_state193_102_2 + shifted_state193_102_4 + shifted_state193_104_0 + shifted_state193_104_1 + shifted_state193_104_2 + shifted_state193_104_4 + shifted_state193_104_6 + shifted_state193_107_3 + shifted_state193_107_4 + shifted_state193_107_5 + shifted_state193_107_6 + shifted_state193_107_7 + shifted_state193_108_0 + shifted_state193_108_2 + shifted_state193_108_5 + shifted_state193_108_6 + shifted_state193_108_7 + shifted_state193_113_0 + shifted_state193_113_1 + shifted_state193_113_5 + shifted_state193_128_0 + shifted_state193_128_1 + shifted_state193_128_4 + shifted_state193_128_5 + shifted_state193_128_6 + shifted_state193_128_7 + shifted_state193_132_1 + shifted_state193_132_3 + shifted_state193_132_5 + shifted_state193_132_6 + shifted_state193_132_7 + shifted_state193_145_0 + shifted_state193_145_1 + shifted_state193_145_3 + shifted_state193_145_4 + shifted_state193_145_5 + shifted_state193_145_6 + shifted_state193_145_7 + shifted_state193_162_1 + shifted_state193_162_3 + shifted_state193_162_4 + shifted_state193_162_6 + shifted_state193_162_7 + shifted_state193_163_0 + shifted_state193_163_2 + shifted_state193_163_5 + shifted_state193_168_0 + shifted_state193_168_1 + shifted_state193_168_4 + shifted_state193_168_5 + shifted_state193_168_6 + shifted_state193_168_7 + shifted_state193_181_2 + shifted_state193_184_3 + shifted_state193_184_5);
      reservoir_sum_parallel[194] = (shifted_state194_10_1 + shifted_state194_10_2 + shifted_state194_10_4 + shifted_state194_30_0 + shifted_state194_30_3 + shifted_state194_30_5 + shifted_state194_31_0 + shifted_state194_31_1 + shifted_state194_31_2 + shifted_state194_31_4 + shifted_state194_31_5 + shifted_state194_31_6 + shifted_state194_31_7 + shifted_state194_32_2 + shifted_state194_32_4 + shifted_state194_122_4 + shifted_state194_122_5 + shifted_state194_127_0 + shifted_state194_127_1 + shifted_state194_127_2 + shifted_state194_127_3 + shifted_state194_127_4 + shifted_state194_127_5 + shifted_state194_127_6 + shifted_state194_127_7 + shifted_state194_155_0 + shifted_state194_155_3 + shifted_state194_155_4 + shifted_state194_155_5 + shifted_state194_155_6 + shifted_state194_155_7 + shifted_state194_179_0 + shifted_state194_179_1 + shifted_state194_179_4 + shifted_state194_179_5 + shifted_state194_179_6 + shifted_state194_179_7 + shifted_state194_183_0 + shifted_state194_183_1 + shifted_state194_183_2 + shifted_state194_189_1 + shifted_state194_189_2 + shifted_state194_189_3 + shifted_state194_189_4 + shifted_state194_189_5 + shifted_state194_189_6 + shifted_state194_189_7);
      reservoir_sum_parallel[195] = (shifted_state195_14_0 + shifted_state195_14_1 + shifted_state195_14_2 + shifted_state195_14_3 + shifted_state195_14_5 + shifted_state195_14_7 + shifted_state195_19_3 + shifted_state195_19_4 + shifted_state195_63_1 + shifted_state195_63_2 + shifted_state195_63_3 + shifted_state195_63_4 + shifted_state195_67_0 + shifted_state195_67_3 + shifted_state195_67_6 + shifted_state195_67_7 + shifted_state195_74_0 + shifted_state195_74_1 + shifted_state195_96_3 + shifted_state195_96_5 + shifted_state195_96_6 + shifted_state195_96_7 + shifted_state195_98_0 + shifted_state195_98_1 + shifted_state195_109_1 + shifted_state195_109_2 + shifted_state195_109_4 + shifted_state195_109_5 + shifted_state195_109_6 + shifted_state195_109_7 + shifted_state195_126_2 + shifted_state195_126_4 + shifted_state195_126_5 + shifted_state195_126_6 + shifted_state195_126_7 + shifted_state195_139_0 + shifted_state195_139_4 + shifted_state195_141_0 + shifted_state195_141_1 + shifted_state195_141_2 + shifted_state195_141_4 + shifted_state195_145_0 + shifted_state195_145_1 + shifted_state195_145_2 + shifted_state195_145_4 + shifted_state195_145_5 + shifted_state195_145_6 + shifted_state195_145_7 + shifted_state195_163_0 + shifted_state195_163_2 + shifted_state195_163_3 + shifted_state195_163_4 + shifted_state195_163_5 + shifted_state195_163_6 + shifted_state195_163_7 + shifted_state195_171_1 + shifted_state195_171_2 + shifted_state195_171_4 + shifted_state195_178_0 + shifted_state195_178_1 + shifted_state195_178_5 + shifted_state195_178_6 + shifted_state195_178_7 + shifted_state195_190_1 + shifted_state195_190_3 + shifted_state195_190_4 + shifted_state195_190_5 + shifted_state195_190_6 + shifted_state195_190_7 + shifted_state195_195_2 + shifted_state195_195_3 + shifted_state195_195_5 + shifted_state195_195_6 + shifted_state195_195_7);
      reservoir_sum_parallel[196] = (shifted_state196_4_0 + shifted_state196_4_2 + shifted_state196_4_3 + shifted_state196_4_4 + shifted_state196_4_5 + shifted_state196_4_6 + shifted_state196_4_7 + shifted_state196_7_1 + shifted_state196_7_4 + shifted_state196_7_5 + shifted_state196_7_6 + shifted_state196_7_7 + shifted_state196_43_1 + shifted_state196_43_4 + shifted_state196_49_0 + shifted_state196_49_2 + shifted_state196_49_3 + shifted_state196_49_5 + shifted_state196_51_1 + shifted_state196_51_2 + shifted_state196_51_3 + shifted_state196_51_4 + shifted_state196_51_5 + shifted_state196_51_6 + shifted_state196_51_7 + shifted_state196_74_0 + shifted_state196_74_4 + shifted_state196_74_5 + shifted_state196_74_6 + shifted_state196_74_7 + shifted_state196_76_1 + shifted_state196_76_5 + shifted_state196_102_1 + shifted_state196_102_4 + shifted_state196_112_0 + shifted_state196_112_1 + shifted_state196_112_2 + shifted_state196_126_0 + shifted_state196_126_2 + shifted_state196_126_4 + shifted_state196_126_5 + shifted_state196_142_1 + shifted_state196_142_2 + shifted_state196_142_4 + shifted_state196_142_5 + shifted_state196_142_6 + shifted_state196_142_7 + shifted_state196_165_0 + shifted_state196_165_1 + shifted_state196_165_3 + shifted_state196_172_0 + shifted_state196_172_3 + shifted_state196_172_4 + shifted_state196_172_6 + shifted_state196_180_0 + shifted_state196_180_1 + shifted_state196_180_2 + shifted_state196_180_3 + shifted_state196_182_1 + shifted_state196_182_4 + shifted_state196_182_5 + shifted_state196_182_6 + shifted_state196_182_7 + shifted_state196_198_3 + shifted_state196_198_4 + shifted_state196_198_6 + shifted_state196_198_7);
      reservoir_sum_parallel[197] = (shifted_state197_0_0 + shifted_state197_0_1 + shifted_state197_0_4 + shifted_state197_0_5 + shifted_state197_0_6 + shifted_state197_0_7 + shifted_state197_44_4 + shifted_state197_87_0 + shifted_state197_87_2 + shifted_state197_87_5 + shifted_state197_89_1 + shifted_state197_89_3 + shifted_state197_89_4 + shifted_state197_89_5 + shifted_state197_89_6 + shifted_state197_89_7 + shifted_state197_90_0 + shifted_state197_90_3 + shifted_state197_90_5 + shifted_state197_121_0 + shifted_state197_121_1 + shifted_state197_121_3 + shifted_state197_121_4 + shifted_state197_121_5 + shifted_state197_121_6 + shifted_state197_121_7 + shifted_state197_137_2 + shifted_state197_137_3 + shifted_state197_137_4 + shifted_state197_137_5 + shifted_state197_137_6 + shifted_state197_137_7 + shifted_state197_141_1 + shifted_state197_141_3 + shifted_state197_141_4 + shifted_state197_141_5 + shifted_state197_143_1 + shifted_state197_143_3 + shifted_state197_143_4 + shifted_state197_143_5 + shifted_state197_143_6 + shifted_state197_143_7 + shifted_state197_150_0 + shifted_state197_150_3 + shifted_state197_150_4 + shifted_state197_150_6 + shifted_state197_150_7 + shifted_state197_152_2 + shifted_state197_156_3 + shifted_state197_156_5 + shifted_state197_156_6 + shifted_state197_156_7 + shifted_state197_159_0 + shifted_state197_159_2 + shifted_state197_159_3 + shifted_state197_159_4 + shifted_state197_159_6 + shifted_state197_159_7 + shifted_state197_163_0 + shifted_state197_163_1 + shifted_state197_163_2 + shifted_state197_163_4 + shifted_state197_163_5 + shifted_state197_176_1 + shifted_state197_176_2 + shifted_state197_176_3 + shifted_state197_195_1 + shifted_state197_195_3 + shifted_state197_195_5 + shifted_state197_195_6 + shifted_state197_195_7);
      reservoir_sum_parallel[198] = (shifted_state198_5_0 + shifted_state198_5_1 + shifted_state198_5_3 + shifted_state198_5_4 + shifted_state198_5_6 + shifted_state198_5_7 + shifted_state198_7_0 + shifted_state198_7_1 + shifted_state198_7_2 + shifted_state198_7_3 + shifted_state198_7_4 + shifted_state198_9_4 + shifted_state198_10_0 + shifted_state198_10_1 + shifted_state198_10_2 + shifted_state198_10_3 + shifted_state198_10_4 + shifted_state198_10_5 + shifted_state198_10_6 + shifted_state198_10_7 + shifted_state198_11_1 + shifted_state198_11_2 + shifted_state198_11_3 + shifted_state198_11_4 + shifted_state198_24_0 + shifted_state198_24_2 + shifted_state198_24_4 + shifted_state198_42_0 + shifted_state198_42_2 + shifted_state198_42_4 + shifted_state198_83_1 + shifted_state198_83_2 + shifted_state198_83_3 + shifted_state198_83_6 + shifted_state198_83_7 + shifted_state198_84_0 + shifted_state198_84_1 + shifted_state198_84_5 + shifted_state198_84_6 + shifted_state198_84_7 + shifted_state198_105_3 + shifted_state198_105_4 + shifted_state198_105_5 + shifted_state198_105_6 + shifted_state198_105_7 + shifted_state198_116_1 + shifted_state198_116_2 + shifted_state198_116_3 + shifted_state198_116_4 + shifted_state198_116_5 + shifted_state198_116_6 + shifted_state198_116_7 + shifted_state198_128_1 + shifted_state198_152_1 + shifted_state198_152_4 + shifted_state198_158_1 + shifted_state198_158_2 + shifted_state198_158_3 + shifted_state198_158_4 + shifted_state198_158_5 + shifted_state198_158_6 + shifted_state198_158_7 + shifted_state198_160_1 + shifted_state198_160_3 + shifted_state198_160_5 + shifted_state198_160_6 + shifted_state198_160_7 + shifted_state198_161_1 + shifted_state198_161_3 + shifted_state198_161_4 + shifted_state198_161_5 + shifted_state198_161_6 + shifted_state198_161_7 + shifted_state198_179_0 + shifted_state198_179_1 + shifted_state198_179_3 + shifted_state198_179_5 + shifted_state198_179_6 + shifted_state198_179_7 + shifted_state198_188_1 + shifted_state198_188_2 + shifted_state198_188_3 + shifted_state198_188_4 + shifted_state198_188_5 + shifted_state198_188_6 + shifted_state198_188_7 + shifted_state198_189_1 + shifted_state198_189_2 + shifted_state198_189_3 + shifted_state198_189_4);
      reservoir_sum_parallel[199] = (shifted_state199_2_1 + shifted_state199_2_4 + shifted_state199_6_0 + shifted_state199_6_1 + shifted_state199_6_2 + shifted_state199_6_5 + shifted_state199_41_0 + shifted_state199_41_2 + shifted_state199_41_4 + shifted_state199_41_6 + shifted_state199_41_7 + shifted_state199_53_1 + shifted_state199_53_3 + shifted_state199_59_1 + shifted_state199_59_2 + shifted_state199_59_4 + shifted_state199_59_6 + shifted_state199_59_7 + shifted_state199_64_0 + shifted_state199_64_1 + shifted_state199_65_1 + shifted_state199_65_2 + shifted_state199_65_4 + shifted_state199_78_0 + shifted_state199_82_2 + shifted_state199_82_4 + shifted_state199_82_6 + shifted_state199_82_7 + shifted_state199_136_0 + shifted_state199_136_4 + shifted_state199_136_5 + shifted_state199_145_0 + shifted_state199_145_1 + shifted_state199_145_3 + shifted_state199_145_4 + shifted_state199_145_5 + shifted_state199_146_0 + shifted_state199_146_2 + shifted_state199_146_3 + shifted_state199_159_2 + shifted_state199_159_3 + shifted_state199_159_4 + shifted_state199_159_5 + shifted_state199_159_6 + shifted_state199_159_7 + shifted_state199_176_1 + shifted_state199_176_2 + shifted_state199_176_4 + shifted_state199_186_1 + shifted_state199_186_2 + shifted_state199_186_3 + shifted_state199_186_4 + shifted_state199_186_5 + shifted_state199_186_6 + shifted_state199_186_7 + shifted_state199_191_1 + shifted_state199_191_5 + shifted_state199_191_6 + shifted_state199_191_7);
      // Threshold comparisons
      for (i = 0; i < num_reservoir_neurons; i = i + 1) begin
          reg_input[i] = 0;
          if (input_sum_parallel[i] < a_scaled) begin
              reg_input[i] = a_scaled;
         end
          else if (input_sum_parallel[i] > b_scaled) begin
              reg_input[i] = b_scaled;
          end
          else begin
              reg_input[i] = input_sum_parallel[i];
          end
      end

      for (k = 0; k < num_reservoir_neurons; k = k + 1) begin
          reg_reservoir[k] = 0;
          if (reservoir_sum_parallel[k] < c_scaled) begin
              reg_reservoir[i] = c_scaled;
          end
          else if (reservoir_sum_parallel[k] > d_scaled) begin
              reg_reservoir[k] = d_scaled;
          end
          else begin
              reg_reservoir[k] = reservoir_sum_parallel[k];
          end
      end


      for (j = 0; j < num_reservoir_neurons; j = j + 1) begin
      reg_input[j]=reg_input[j]+16'd1628;

          reg_input[j] = reg_input[j] >> 8;
          reg_reservoir[j]=reg_reservoir[j]+16'd17641;
          reg_reservoir[j]= reg_reservoir[j] >> 8;
      end

  // Store results in reservoir_states
      for (m = 0; m < num_reservoir_neurons; m = m + 1) begin
          reservoir_state[m] <= reg_reservoir[m] + reg_input[m]-255;
      end
      // Output calculation
      output_sum = 0;
      output_sum = output_sum + (shifted_state_out0_0 + shifted_state_out0_2 + shifted_state_out0_3 + shifted_state_out0_4 + shifted_state_out0_5 + shifted_state_out0_6 + shifted_state_out0_7 + shifted_state_out1_0 + shifted_state_out1_2 + shifted_state_out2_2 + shifted_state_out3_1 + shifted_state_out5_1 + shifted_state_out5_2 + shifted_state_out5_3 + shifted_state_out5_4 + shifted_state_out5_5 + shifted_state_out5_6 + shifted_state_out5_7 + shifted_state_out6_1 + shifted_state_out7_1 + shifted_state_out7_3 + shifted_state_out7_4 + shifted_state_out7_5 + shifted_state_out7_6 + shifted_state_out7_7 + shifted_state_out9_2 + shifted_state_out10_1 + shifted_state_out11_0 + shifted_state_out11_2 + shifted_state_out12_1 + shifted_state_out13_0 + shifted_state_out13_2 + shifted_state_out13_3 + shifted_state_out13_4 + shifted_state_out13_5 + shifted_state_out13_6 + shifted_state_out13_7 + shifted_state_out14_0 + shifted_state_out14_1 + shifted_state_out15_0 + shifted_state_out15_4 + shifted_state_out16_0 + shifted_state_out16_2 + shifted_state_out16_4 + shifted_state_out16_5 + shifted_state_out16_6 + shifted_state_out16_7 + shifted_state_out17_1 + shifted_state_out17_2 + shifted_state_out17_3 + shifted_state_out17_4 + shifted_state_out17_5 + shifted_state_out17_6 + shifted_state_out17_7 + shifted_state_out18_0 + shifted_state_out18_1 + shifted_state_out19_0 + shifted_state_out19_1 + shifted_state_out19_2 + shifted_state_out19_3 + shifted_state_out20_2 + shifted_state_out21_0 + shifted_state_out21_1 + shifted_state_out21_2 + shifted_state_out21_3 + shifted_state_out21_4 + shifted_state_out21_5 + shifted_state_out21_6 + shifted_state_out21_7 + shifted_state_out22_0 + shifted_state_out22_1 + shifted_state_out23_3 + shifted_state_out24_1 + shifted_state_out25_1 + shifted_state_out25_4 + shifted_state_out25_5 + shifted_state_out26_1 + shifted_state_out26_2 + shifted_state_out27_1 + shifted_state_out27_2 + shifted_state_out28_0 + shifted_state_out28_2 + shifted_state_out30_1 + shifted_state_out30_2 + shifted_state_out30_3 + shifted_state_out30_4 + shifted_state_out30_5 + shifted_state_out30_6 + shifted_state_out30_7 + shifted_state_out31_3 + shifted_state_out32_0 + shifted_state_out32_1 + shifted_state_out32_3 + shifted_state_out32_4 + shifted_state_out32_5 + shifted_state_out32_6 + shifted_state_out32_7 + shifted_state_out33_1 + shifted_state_out34_2 + shifted_state_out35_0 + shifted_state_out35_1 + shifted_state_out35_2 + shifted_state_out36_1 + shifted_state_out36_2 + shifted_state_out36_3 + shifted_state_out36_4 + shifted_state_out36_5 + shifted_state_out36_6 + shifted_state_out36_7 + shifted_state_out37_0 + shifted_state_out37_1 + shifted_state_out38_1 + shifted_state_out38_3 + shifted_state_out38_4 + shifted_state_out38_5 + shifted_state_out38_6 + shifted_state_out38_7 + shifted_state_out39_1 + shifted_state_out39_3 + shifted_state_out39_4 + shifted_state_out39_5 + shifted_state_out39_6 + shifted_state_out39_7 + shifted_state_out40_1 + shifted_state_out42_0 + shifted_state_out42_3 + shifted_state_out43_0 + shifted_state_out43_1 + shifted_state_out43_2 + shifted_state_out43_3 + shifted_state_out43_4 + shifted_state_out43_5 + shifted_state_out43_6 + shifted_state_out43_7 + shifted_state_out44_1 + shifted_state_out45_2 + shifted_state_out45_3 + shifted_state_out45_4 + shifted_state_out45_5 + shifted_state_out45_6 + shifted_state_out45_7 + shifted_state_out46_0 + shifted_state_out46_3 + shifted_state_out46_4 + shifted_state_out46_5 + shifted_state_out46_6 + shifted_state_out46_7 + shifted_state_out47_0 + shifted_state_out47_1 + shifted_state_out48_1 + shifted_state_out48_2 + shifted_state_out48_3 + shifted_state_out48_4 + shifted_state_out48_5 + shifted_state_out48_6 + shifted_state_out48_7 + shifted_state_out50_1 + shifted_state_out50_2 + shifted_state_out51_0 + shifted_state_out51_3 + shifted_state_out52_0 + shifted_state_out52_2 + shifted_state_out52_3 + shifted_state_out52_4 + shifted_state_out52_5 + shifted_state_out52_6 + shifted_state_out52_7 + shifted_state_out53_0 + shifted_state_out53_1 + shifted_state_out53_2 + shifted_state_out55_0 + shifted_state_out55_1 + shifted_state_out55_3 + shifted_state_out55_4 + shifted_state_out55_5 + shifted_state_out55_6 + shifted_state_out55_7 + shifted_state_out56_1 + shifted_state_out57_0 + shifted_state_out57_1 + shifted_state_out57_2 + shifted_state_out58_0 + shifted_state_out58_2 + shifted_state_out58_3 + shifted_state_out58_4 + shifted_state_out58_5 + shifted_state_out58_6 + shifted_state_out58_7 + shifted_state_out59_0 + shifted_state_out59_1 + shifted_state_out61_0 + shifted_state_out62_1 + shifted_state_out62_2 + shifted_state_out62_3 + shifted_state_out62_4 + shifted_state_out62_5 + shifted_state_out62_6 + shifted_state_out62_7 + shifted_state_out63_3 + shifted_state_out64_1 + shifted_state_out64_2 + shifted_state_out64_3 + shifted_state_out64_4 + shifted_state_out64_5 + shifted_state_out64_6 + shifted_state_out64_7 + shifted_state_out65_0 + shifted_state_out65_2 + shifted_state_out66_1 + shifted_state_out67_0 + shifted_state_out69_0 + shifted_state_out70_1 + shifted_state_out70_3 + shifted_state_out70_4 + shifted_state_out70_5 + shifted_state_out70_6 + shifted_state_out70_7 + shifted_state_out71_1 + shifted_state_out72_0 + shifted_state_out72_1 + shifted_state_out72_3 + shifted_state_out72_4 + shifted_state_out72_5 + shifted_state_out72_6 + shifted_state_out72_7 + shifted_state_out73_0 + shifted_state_out73_1 + shifted_state_out73_3 + shifted_state_out73_4 + shifted_state_out73_5 + shifted_state_out73_6 + shifted_state_out73_7 + shifted_state_out74_0 + shifted_state_out74_2 + shifted_state_out75_0 + shifted_state_out76_1 + shifted_state_out76_2 + shifted_state_out76_3 + shifted_state_out76_4 + shifted_state_out76_5 + shifted_state_out76_6 + shifted_state_out76_7 + shifted_state_out77_2 + shifted_state_out77_3 + shifted_state_out77_4 + shifted_state_out77_5 + shifted_state_out77_6 + shifted_state_out77_7 + shifted_state_out78_0 + shifted_state_out78_1 + shifted_state_out78_2 + shifted_state_out78_3 + shifted_state_out78_4 + shifted_state_out78_5 + shifted_state_out78_6 + shifted_state_out78_7 + shifted_state_out79_1 + shifted_state_out79_2 + shifted_state_out79_3 + shifted_state_out79_4 + shifted_state_out79_5 + shifted_state_out79_6 + shifted_state_out79_7 + shifted_state_out80_0 + shifted_state_out80_1 + shifted_state_out80_2 + shifted_state_out81_0 + shifted_state_out82_0 + shifted_state_out82_1 + shifted_state_out82_2 + shifted_state_out82_3 + shifted_state_out82_4 + shifted_state_out82_5 + shifted_state_out82_6 + shifted_state_out82_7 + shifted_state_out83_2 + shifted_state_out83_3 + shifted_state_out83_4 + shifted_state_out83_5 + shifted_state_out83_6 + shifted_state_out83_7 + shifted_state_out84_3 + shifted_state_out84_4 + shifted_state_out84_5 + shifted_state_out84_6 + shifted_state_out84_7 + shifted_state_out85_0 + shifted_state_out86_2 + shifted_state_out87_3 + shifted_state_out87_4 + shifted_state_out87_5 + shifted_state_out87_6 + shifted_state_out87_7 + shifted_state_out88_0 + shifted_state_out89_2 + shifted_state_out89_3 + shifted_state_out90_3 + shifted_state_out91_0 + shifted_state_out91_1 + shifted_state_out91_3 + shifted_state_out91_4 + shifted_state_out91_5 + shifted_state_out91_6 + shifted_state_out91_7 + shifted_state_out92_0 + shifted_state_out92_2 + shifted_state_out93_0 + shifted_state_out93_1 + shifted_state_out93_2 + shifted_state_out93_3 + shifted_state_out93_4 + shifted_state_out93_5 + shifted_state_out93_6 + shifted_state_out93_7 + shifted_state_out95_0 + shifted_state_out95_1 + shifted_state_out95_2 + shifted_state_out95_3 + shifted_state_out95_4 + shifted_state_out95_5 + shifted_state_out95_6 + shifted_state_out95_7 + shifted_state_out96_0 + shifted_state_out96_2 + shifted_state_out97_0 + shifted_state_out97_1 + shifted_state_out97_2 + shifted_state_out97_3 + shifted_state_out97_4 + shifted_state_out97_5 + shifted_state_out97_6 + shifted_state_out97_7 + shifted_state_out98_2 + shifted_state_out100_0 + shifted_state_out100_1 + shifted_state_out100_3 + shifted_state_out100_4 + shifted_state_out100_5 + shifted_state_out100_6 + shifted_state_out100_7 + shifted_state_out101_1 + shifted_state_out102_1 + shifted_state_out102_2 + shifted_state_out102_3 + shifted_state_out102_4 + shifted_state_out102_5 + shifted_state_out102_6 + shifted_state_out102_7 + shifted_state_out103_1 + shifted_state_out103_2 + shifted_state_out103_3 + shifted_state_out103_4 + shifted_state_out103_5 + shifted_state_out103_6 + shifted_state_out103_7 + shifted_state_out105_0 + shifted_state_out105_2 + shifted_state_out106_0 + shifted_state_out106_1 + shifted_state_out107_0 + shifted_state_out108_0 + shifted_state_out108_3 + shifted_state_out109_2 + shifted_state_out109_3 + shifted_state_out109_4 + shifted_state_out109_5 + shifted_state_out109_6 + shifted_state_out109_7 + shifted_state_out111_0 + shifted_state_out111_1 + shifted_state_out112_1 + shifted_state_out112_3 + shifted_state_out112_4 + shifted_state_out112_5 + shifted_state_out112_6 + shifted_state_out112_7 + shifted_state_out113_1 + shifted_state_out113_3 + shifted_state_out113_4 + shifted_state_out113_5 + shifted_state_out113_6 + shifted_state_out113_7 + shifted_state_out114_0 + shifted_state_out114_2 + shifted_state_out114_3 + shifted_state_out114_4 + shifted_state_out114_5 + shifted_state_out114_6 + shifted_state_out114_7 + shifted_state_out115_1 + shifted_state_out115_3 + shifted_state_out115_4 + shifted_state_out115_5 + shifted_state_out115_6 + shifted_state_out115_7 + shifted_state_out116_0 + shifted_state_out117_0 + shifted_state_out117_2 + shifted_state_out118_1 + shifted_state_out118_2 + shifted_state_out119_0 + shifted_state_out119_1 + shifted_state_out119_2 + shifted_state_out119_3 + shifted_state_out119_4 + shifted_state_out119_5 + shifted_state_out119_6 + shifted_state_out119_7 + shifted_state_out120_0 + shifted_state_out120_1 + shifted_state_out120_3 + shifted_state_out120_4 + shifted_state_out120_5 + shifted_state_out120_6 + shifted_state_out120_7 + shifted_state_out121_0 + shifted_state_out121_2 + shifted_state_out121_3 + shifted_state_out121_4 + shifted_state_out121_5 + shifted_state_out121_6 + shifted_state_out121_7 + shifted_state_out122_0 + shifted_state_out122_2 + shifted_state_out123_0 + shifted_state_out123_1 + shifted_state_out124_1 + shifted_state_out124_2 + shifted_state_out124_3 + shifted_state_out124_4 + shifted_state_out124_5 + shifted_state_out124_6 + shifted_state_out124_7 + shifted_state_out125_0 + shifted_state_out125_1 + shifted_state_out125_2 + shifted_state_out125_3 + shifted_state_out125_4 + shifted_state_out125_5 + shifted_state_out125_6 + shifted_state_out125_7 + shifted_state_out126_1 + shifted_state_out126_2 + shifted_state_out127_1 + shifted_state_out128_0 + shifted_state_out128_1 + shifted_state_out129_1 + shifted_state_out129_2 + shifted_state_out129_3 + shifted_state_out129_4 + shifted_state_out129_5 + shifted_state_out129_6 + shifted_state_out129_7 + shifted_state_out131_0 + shifted_state_out132_0 + shifted_state_out133_0 + shifted_state_out133_1 + shifted_state_out134_1 + shifted_state_out134_2 + shifted_state_out135_0 + shifted_state_out135_1 + shifted_state_out135_2 + shifted_state_out135_3 + shifted_state_out135_4 + shifted_state_out135_5 + shifted_state_out135_6 + shifted_state_out135_7 + shifted_state_out137_0 + shifted_state_out137_2 + shifted_state_out138_2 + shifted_state_out138_3 + shifted_state_out138_4 + shifted_state_out138_5 + shifted_state_out138_6 + shifted_state_out138_7 + shifted_state_out139_0 + shifted_state_out139_1 + shifted_state_out139_2 + shifted_state_out139_3 + shifted_state_out139_4 + shifted_state_out139_5 + shifted_state_out139_6 + shifted_state_out139_7 + shifted_state_out140_0 + shifted_state_out140_1 + shifted_state_out140_2 + shifted_state_out140_3 + shifted_state_out140_4 + shifted_state_out140_5 + shifted_state_out140_6 + shifted_state_out140_7 + shifted_state_out141_2 + shifted_state_out142_1 + shifted_state_out142_2 + shifted_state_out142_3 + shifted_state_out142_4 + shifted_state_out142_5 + shifted_state_out142_6 + shifted_state_out142_7 + shifted_state_out143_0 + shifted_state_out143_1 + shifted_state_out143_2 + shifted_state_out143_3 + shifted_state_out143_4 + shifted_state_out143_5 + shifted_state_out143_6 + shifted_state_out143_7 + shifted_state_out144_2 + shifted_state_out144_3 + shifted_state_out144_4 + shifted_state_out144_5 + shifted_state_out144_6 + shifted_state_out144_7 + shifted_state_out145_0 + shifted_state_out145_1 + shifted_state_out145_2 + shifted_state_out145_3 + shifted_state_out145_4 + shifted_state_out145_5 + shifted_state_out145_6 + shifted_state_out145_7 + shifted_state_out146_0 + shifted_state_out146_1 + shifted_state_out146_3 + shifted_state_out146_4 + shifted_state_out146_5 + shifted_state_out146_6 + shifted_state_out146_7 + shifted_state_out147_0 + shifted_state_out147_1 + shifted_state_out147_2 + shifted_state_out148_1 + shifted_state_out149_1 + shifted_state_out149_3 + shifted_state_out150_0 + shifted_state_out150_2 + shifted_state_out150_3 + shifted_state_out150_4 + shifted_state_out150_5 + shifted_state_out150_6 + shifted_state_out150_7 + shifted_state_out151_1 + shifted_state_out151_2 + shifted_state_out151_3 + shifted_state_out151_4 + shifted_state_out151_5 + shifted_state_out151_6 + shifted_state_out151_7 + shifted_state_out152_1 + shifted_state_out152_2 + shifted_state_out152_3 + shifted_state_out152_4 + shifted_state_out152_5 + shifted_state_out152_6 + shifted_state_out152_7 + shifted_state_out153_0 + shifted_state_out153_2 + shifted_state_out153_3 + shifted_state_out153_4 + shifted_state_out153_5 + shifted_state_out153_6 + shifted_state_out153_7 + shifted_state_out154_1 + shifted_state_out154_2 + shifted_state_out154_3 + shifted_state_out154_4 + shifted_state_out154_5 + shifted_state_out154_6 + shifted_state_out154_7 + shifted_state_out155_0 + shifted_state_out155_7 + shifted_state_out156_3 + shifted_state_out156_4 + shifted_state_out156_5 + shifted_state_out156_6 + shifted_state_out156_7 + shifted_state_out157_1 + shifted_state_out157_2 + shifted_state_out157_3 + shifted_state_out157_4 + shifted_state_out157_5 + shifted_state_out157_6 + shifted_state_out157_7 + shifted_state_out158_2 + shifted_state_out158_3 + shifted_state_out158_4 + shifted_state_out158_5 + shifted_state_out158_6 + shifted_state_out158_7 + shifted_state_out159_0 + shifted_state_out159_2 + shifted_state_out160_2 + shifted_state_out160_3 + shifted_state_out160_4 + shifted_state_out160_5 + shifted_state_out160_6 + shifted_state_out160_7 + shifted_state_out161_0 + shifted_state_out161_1 + shifted_state_out161_2 + shifted_state_out161_3 + shifted_state_out161_4 + shifted_state_out161_5 + shifted_state_out161_6 + shifted_state_out161_7 + shifted_state_out162_1 + shifted_state_out162_2 + shifted_state_out162_3 + shifted_state_out162_4 + shifted_state_out162_5 + shifted_state_out162_6 + shifted_state_out162_7 + shifted_state_out164_0 + shifted_state_out164_3 + shifted_state_out164_4 + shifted_state_out164_5 + shifted_state_out164_6 + shifted_state_out164_7 + shifted_state_out165_0 + shifted_state_out165_2 + shifted_state_out166_0 + shifted_state_out166_1 + shifted_state_out166_3 + shifted_state_out166_4 + shifted_state_out166_5 + shifted_state_out166_6 + shifted_state_out166_7 + shifted_state_out167_1 + shifted_state_out167_2 + shifted_state_out167_3 + shifted_state_out167_4 + shifted_state_out167_5 + shifted_state_out167_6 + shifted_state_out167_7 + shifted_state_out169_1 + shifted_state_out170_0 + shifted_state_out170_2 + shifted_state_out171_2 + shifted_state_out172_1 + shifted_state_out173_1 + shifted_state_out173_2 + shifted_state_out174_3 + shifted_state_out174_4 + shifted_state_out174_5 + shifted_state_out174_6 + shifted_state_out174_7 + shifted_state_out175_0 + shifted_state_out175_1 + shifted_state_out176_0 + shifted_state_out176_1 + shifted_state_out177_1 + shifted_state_out177_2 + shifted_state_out178_0 + shifted_state_out178_2 + shifted_state_out178_4 + shifted_state_out178_5 + shifted_state_out178_6 + shifted_state_out178_7 + shifted_state_out179_3 + shifted_state_out179_4 + shifted_state_out179_5 + shifted_state_out179_6 + shifted_state_out179_7 + shifted_state_out180_0 + shifted_state_out180_1 + shifted_state_out181_3 + shifted_state_out181_4 + shifted_state_out181_5 + shifted_state_out181_6 + shifted_state_out181_7 + shifted_state_out182_0 + shifted_state_out182_3 + shifted_state_out183_0 + shifted_state_out183_2 + shifted_state_out183_3 + shifted_state_out183_4 + shifted_state_out183_5 + shifted_state_out183_6 + shifted_state_out183_7 + shifted_state_out184_0 + shifted_state_out184_1 + shifted_state_out185_0 + shifted_state_out185_1 + shifted_state_out185_2 + shifted_state_out186_2 + shifted_state_out186_3 + shifted_state_out186_4 + shifted_state_out186_5 + shifted_state_out186_6 + shifted_state_out186_7 + shifted_state_out187_1 + shifted_state_out188_0 + shifted_state_out188_2 + shifted_state_out188_3 + shifted_state_out188_4 + shifted_state_out188_5 + shifted_state_out188_6 + shifted_state_out188_7 + shifted_state_out189_1 + shifted_state_out190_1 + shifted_state_out190_2 + shifted_state_out190_3 + shifted_state_out190_4 + shifted_state_out190_5 + shifted_state_out190_6 + shifted_state_out190_7 + shifted_state_out191_1 + shifted_state_out192_0 + shifted_state_out193_0 + shifted_state_out193_2 + shifted_state_out193_3 + shifted_state_out193_4 + shifted_state_out193_5 + shifted_state_out193_6 + shifted_state_out193_7 + shifted_state_out194_0 + shifted_state_out194_1 + shifted_state_out194_2 + shifted_state_out194_3 + shifted_state_out194_4 + shifted_state_out194_5 + shifted_state_out194_6 + shifted_state_out194_7 + shifted_state_out195_0 + shifted_state_out195_1 + shifted_state_out195_2 + shifted_state_out195_3 + shifted_state_out195_4 + shifted_state_out195_5 + shifted_state_out195_6 + shifted_state_out195_7 + shifted_state_out196_1 + shifted_state_out196_2 + shifted_state_out196_3 + shifted_state_out196_4 + shifted_state_out196_5 + shifted_state_out196_6 + shifted_state_out196_7 + shifted_state_out197_1 + shifted_state_out197_2 + shifted_state_out197_3 + shifted_state_out197_4 + shifted_state_out197_5 + shifted_state_out197_6 + shifted_state_out197_7 + shifted_state_out198_0 + shifted_state_out198_1 + shifted_state_out198_3 + shifted_state_out198_4 + shifted_state_out198_5 + shifted_state_out198_6 + shifted_state_out198_7 + shifted_state_out199_0 + shifted_state_out199_1 + shifted_state_out199_3 + shifted_state_out199_4 + shifted_state_out199_5 + shifted_state_out199_6 + shifted_state_out199_7);

    end
    assign output_data = output_sum;
endmodule
